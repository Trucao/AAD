module jogo(
	input advance_clk,
	input reset,
	input [5:0] row,
	input [5:0] column,
	output pixel
);
	parameter ROWS = 48;
	parameter COLUMNS = 64;

	reg [COLUMNS-1:0] board [0:ROWS-1];
	reg [COLUMNS-1:0] next_board [0:ROWS-1];
	
	always @(posedge advance_clk or posedge reset) begin
		integer i, j;
	
		if (reset) begin
		   board[0][0] <= 0;
		   board[0][1] <= 0;
		   board[0][2] <= 0;
		   board[0][3] <= 0;
		   board[0][4] <= 0;
		   board[0][5] <= 0;
		   board[0][6] <= 0;
		   board[0][7] <= 0;
		   board[0][8] <= 0;
		   board[0][9] <= 0;
		   board[0][10] <= 0;
		   board[0][11] <= 0;
		   board[0][12] <= 0;
		   board[0][13] <= 0;
		   board[0][14] <= 0;
		   board[0][15] <= 0;
		   board[0][16] <= 0;
		   board[0][17] <= 0;
		   board[0][18] <= 0;
		   board[0][19] <= 0;
		   board[0][20] <= 0;
		   board[0][21] <= 0;
		   board[0][22] <= 0;
		   board[0][23] <= 0;
		   board[0][24] <= 0;
		   board[0][25] <= 0;
		   board[0][26] <= 0;
		   board[0][27] <= 0;
		   board[0][28] <= 0;
		   board[0][29] <= 0;
		   board[0][30] <= 0;
		   board[0][31] <= 0;
		   board[0][32] <= 0;
		   board[0][33] <= 0;
		   board[0][34] <= 0;
		   board[0][35] <= 0;
		   board[0][36] <= 0;
		   board[0][37] <= 0;
		   board[0][38] <= 0;
		   board[0][39] <= 0;
		   board[0][40] <= 0;
		   board[0][41] <= 0;
		   board[0][42] <= 0;
		   board[0][43] <= 0;
		   board[0][44] <= 0;
		   board[0][45] <= 0;
		   board[0][46] <= 0;
		   board[0][47] <= 0;
		   board[0][48] <= 0;
		   board[0][49] <= 0;
		   board[0][50] <= 0;
		   board[0][51] <= 0;
		   board[0][52] <= 0;
		   board[0][53] <= 0;
		   board[0][54] <= 0;
		   board[0][55] <= 0;
		   board[0][56] <= 0;
		   board[0][57] <= 0;
		   board[0][58] <= 0;
		   board[0][59] <= 0;
		   board[0][60] <= 0;
		   board[0][61] <= 0;
		   board[0][62] <= 0;
		   board[0][63] <= 0;
		   board[1][0] <= 0;
		   board[1][1] <= 0;
		   board[1][2] <= 0;
		   board[1][3] <= 0;
		   board[1][4] <= 0;
		   board[1][5] <= 0;
		   board[1][6] <= 0;
		   board[1][7] <= 0;
		   board[1][8] <= 0;
		   board[1][9] <= 0;
		   board[1][10] <= 0;
		   board[1][11] <= 0;
		   board[1][12] <= 0;
		   board[1][13] <= 0;
		   board[1][14] <= 0;
		   board[1][15] <= 0;
		   board[1][16] <= 0;
		   board[1][17] <= 0;
		   board[1][18] <= 0;
		   board[1][19] <= 0;
		   board[1][20] <= 0;
		   board[1][21] <= 0;
		   board[1][22] <= 0;
		   board[1][23] <= 0;
		   board[1][24] <= 0;
		   board[1][25] <= 0;
		   board[1][26] <= 0;
		   board[1][27] <= 0;
		   board[1][28] <= 0;
		   board[1][29] <= 0;
		   board[1][30] <= 0;
		   board[1][31] <= 0;
		   board[1][32] <= 0;
		   board[1][33] <= 0;
		   board[1][34] <= 0;
		   board[1][35] <= 0;
		   board[1][36] <= 0;
		   board[1][37] <= 0;
		   board[1][38] <= 0;
		   board[1][39] <= 0;
		   board[1][40] <= 0;
		   board[1][41] <= 0;
		   board[1][42] <= 0;
		   board[1][43] <= 0;
		   board[1][44] <= 0;
		   board[1][45] <= 0;
		   board[1][46] <= 0;
		   board[1][47] <= 0;
		   board[1][48] <= 0;
		   board[1][49] <= 0;
		   board[1][50] <= 0;
		   board[1][51] <= 0;
		   board[1][52] <= 0;
		   board[1][53] <= 0;
		   board[1][54] <= 0;
		   board[1][55] <= 0;
		   board[1][56] <= 0;
		   board[1][57] <= 0;
		   board[1][58] <= 0;
		   board[1][59] <= 0;
		   board[1][60] <= 0;
		   board[1][61] <= 0;
		   board[1][62] <= 0;
		   board[1][63] <= 0;
		   board[2][0] <= 0;
		   board[2][1] <= 0;
		   board[2][2] <= 0;
		   board[2][3] <= 0;
		   board[2][4] <= 0;
		   board[2][5] <= 0;
		   board[2][6] <= 0;
		   board[2][7] <= 0;
		   board[2][8] <= 0;
		   board[2][9] <= 0;
		   board[2][10] <= 0;
		   board[2][11] <= 0;
		   board[2][12] <= 0;
		   board[2][13] <= 0;
		   board[2][14] <= 0;
		   board[2][15] <= 0;
		   board[2][16] <= 0;
		   board[2][17] <= 0;
		   board[2][18] <= 0;
		   board[2][19] <= 0;
		   board[2][20] <= 0;
		   board[2][21] <= 0;
		   board[2][22] <= 0;
		   board[2][23] <= 0;
		   board[2][24] <= 0;
		   board[2][25] <= 0;
		   board[2][26] <= 0;
		   board[2][27] <= 0;
		   board[2][28] <= 0;
		   board[2][29] <= 0;
		   board[2][30] <= 0;
		   board[2][31] <= 0;
		   board[2][32] <= 0;
		   board[2][33] <= 0;
		   board[2][34] <= 0;
		   board[2][35] <= 0;
		   board[2][36] <= 0;
		   board[2][37] <= 0;
		   board[2][38] <= 0;
		   board[2][39] <= 0;
		   board[2][40] <= 0;
		   board[2][41] <= 0;
		   board[2][42] <= 0;
		   board[2][43] <= 0;
		   board[2][44] <= 0;
		   board[2][45] <= 0;
		   board[2][46] <= 0;
		   board[2][47] <= 0;
		   board[2][48] <= 0;
		   board[2][49] <= 0;
		   board[2][50] <= 0;
		   board[2][51] <= 0;
		   board[2][52] <= 0;
		   board[2][53] <= 0;
		   board[2][54] <= 0;
		   board[2][55] <= 0;
		   board[2][56] <= 0;
		   board[2][57] <= 0;
		   board[2][58] <= 0;
		   board[2][59] <= 0;
		   board[2][60] <= 0;
		   board[2][61] <= 0;
		   board[2][62] <= 0;
		   board[2][63] <= 0;
		   board[3][0] <= 0;
		   board[3][1] <= 0;
		   board[3][2] <= 0;
		   board[3][3] <= 0;
		   board[3][4] <= 0;
		   board[3][5] <= 0;
		   board[3][6] <= 0;
		   board[3][7] <= 0;
		   board[3][8] <= 0;
		   board[3][9] <= 0;
		   board[3][10] <= 0;
		   board[3][11] <= 0;
		   board[3][12] <= 0;
		   board[3][13] <= 0;
		   board[3][14] <= 0;
		   board[3][15] <= 0;
		   board[3][16] <= 0;
		   board[3][17] <= 0;
		   board[3][18] <= 0;
		   board[3][19] <= 0;
		   board[3][20] <= 0;
		   board[3][21] <= 0;
		   board[3][22] <= 0;
		   board[3][23] <= 0;
		   board[3][24] <= 0;
		   board[3][25] <= 0;
		   board[3][26] <= 0;
		   board[3][27] <= 0;
		   board[3][28] <= 0;
		   board[3][29] <= 0;
		   board[3][30] <= 0;
		   board[3][31] <= 0;
		   board[3][32] <= 0;
		   board[3][33] <= 0;
		   board[3][34] <= 0;
		   board[3][35] <= 0;
		   board[3][36] <= 0;
		   board[3][37] <= 0;
		   board[3][38] <= 0;
		   board[3][39] <= 0;
		   board[3][40] <= 0;
		   board[3][41] <= 0;
		   board[3][42] <= 0;
		   board[3][43] <= 0;
		   board[3][44] <= 0;
		   board[3][45] <= 0;
		   board[3][46] <= 0;
		   board[3][47] <= 0;
		   board[3][48] <= 0;
		   board[3][49] <= 0;
		   board[3][50] <= 0;
		   board[3][51] <= 0;
		   board[3][52] <= 0;
		   board[3][53] <= 0;
		   board[3][54] <= 0;
		   board[3][55] <= 0;
		   board[3][56] <= 0;
		   board[3][57] <= 0;
		   board[3][58] <= 0;
		   board[3][59] <= 0;
		   board[3][60] <= 0;
		   board[3][61] <= 0;
		   board[3][62] <= 0;
		   board[3][63] <= 0;
		   board[4][0] <= 0;
		   board[4][1] <= 0;
		   board[4][2] <= 0;
		   board[4][3] <= 0;
		   board[4][4] <= 0;
		   board[4][5] <= 0;
		   board[4][6] <= 0;
		   board[4][7] <= 0;
		   board[4][8] <= 0;
		   board[4][9] <= 0;
		   board[4][10] <= 0;
		   board[4][11] <= 0;
		   board[4][12] <= 0;
		   board[4][13] <= 0;
		   board[4][14] <= 0;
		   board[4][15] <= 0;
		   board[4][16] <= 0;
		   board[4][17] <= 0;
		   board[4][18] <= 0;
		   board[4][19] <= 0;
		   board[4][20] <= 0;
		   board[4][21] <= 0;
		   board[4][22] <= 0;
		   board[4][23] <= 0;
		   board[4][24] <= 0;
		   board[4][25] <= 0;
		   board[4][26] <= 0;
		   board[4][27] <= 0;
		   board[4][28] <= 0;
		   board[4][29] <= 0;
		   board[4][30] <= 0;
		   board[4][31] <= 0;
		   board[4][32] <= 0;
		   board[4][33] <= 0;
		   board[4][34] <= 0;
		   board[4][35] <= 0;
		   board[4][36] <= 0;
		   board[4][37] <= 0;
		   board[4][38] <= 0;
		   board[4][39] <= 0;
		   board[4][40] <= 0;
		   board[4][41] <= 0;
		   board[4][42] <= 0;
		   board[4][43] <= 0;
		   board[4][44] <= 0;
		   board[4][45] <= 0;
		   board[4][46] <= 0;
		   board[4][47] <= 0;
		   board[4][48] <= 0;
		   board[4][49] <= 0;
		   board[4][50] <= 0;
		   board[4][51] <= 0;
		   board[4][52] <= 0;
		   board[4][53] <= 0;
		   board[4][54] <= 0;
		   board[4][55] <= 0;
		   board[4][56] <= 0;
		   board[4][57] <= 0;
		   board[4][58] <= 0;
		   board[4][59] <= 0;
		   board[4][60] <= 0;
		   board[4][61] <= 0;
		   board[4][62] <= 0;
		   board[4][63] <= 0;
		   board[5][0] <= 0;
		   board[5][1] <= 0;
		   board[5][2] <= 0;
		   board[5][3] <= 0;
		   board[5][4] <= 0;
		   board[5][5] <= 0;
		   board[5][6] <= 0;
		   board[5][7] <= 0;
		   board[5][8] <= 0;
		   board[5][9] <= 0;
		   board[5][10] <= 0;
		   board[5][11] <= 0;
		   board[5][12] <= 0;
		   board[5][13] <= 0;
		   board[5][14] <= 0;
		   board[5][15] <= 0;
		   board[5][16] <= 0;
		   board[5][17] <= 0;
		   board[5][18] <= 0;
		   board[5][19] <= 0;
		   board[5][20] <= 0;
		   board[5][21] <= 0;
		   board[5][22] <= 0;
		   board[5][23] <= 0;
		   board[5][24] <= 0;
		   board[5][25] <= 0;
		   board[5][26] <= 0;
		   board[5][27] <= 0;
		   board[5][28] <= 0;
		   board[5][29] <= 0;
		   board[5][30] <= 0;
		   board[5][31] <= 0;
		   board[5][32] <= 0;
		   board[5][33] <= 0;
		   board[5][34] <= 0;
		   board[5][35] <= 0;
		   board[5][36] <= 0;
		   board[5][37] <= 0;
		   board[5][38] <= 0;
		   board[5][39] <= 0;
		   board[5][40] <= 0;
		   board[5][41] <= 0;
		   board[5][42] <= 0;
		   board[5][43] <= 0;
		   board[5][44] <= 0;
		   board[5][45] <= 0;
		   board[5][46] <= 0;
		   board[5][47] <= 0;
		   board[5][48] <= 0;
		   board[5][49] <= 0;
		   board[5][50] <= 0;
		   board[5][51] <= 0;
		   board[5][52] <= 0;
		   board[5][53] <= 0;
		   board[5][54] <= 0;
		   board[5][55] <= 0;
		   board[5][56] <= 0;
		   board[5][57] <= 0;
		   board[5][58] <= 0;
		   board[5][59] <= 0;
		   board[5][60] <= 0;
		   board[5][61] <= 0;
		   board[5][62] <= 0;
		   board[5][63] <= 0;
		   board[6][0] <= 0;
		   board[6][1] <= 0;
		   board[6][2] <= 0;
		   board[6][3] <= 0;
		   board[6][4] <= 0;
		   board[6][5] <= 0;
		   board[6][6] <= 0;
		   board[6][7] <= 0;
		   board[6][8] <= 0;
		   board[6][9] <= 0;
		   board[6][10] <= 0;
		   board[6][11] <= 0;
		   board[6][12] <= 0;
		   board[6][13] <= 0;
		   board[6][14] <= 0;
		   board[6][15] <= 0;
		   board[6][16] <= 0;
		   board[6][17] <= 0;
		   board[6][18] <= 0;
		   board[6][19] <= 0;
		   board[6][20] <= 0;
		   board[6][21] <= 0;
		   board[6][22] <= 0;
		   board[6][23] <= 0;
		   board[6][24] <= 0;
		   board[6][25] <= 0;
		   board[6][26] <= 0;
		   board[6][27] <= 0;
		   board[6][28] <= 0;
		   board[6][29] <= 0;
		   board[6][30] <= 0;
		   board[6][31] <= 0;
		   board[6][32] <= 0;
		   board[6][33] <= 0;
		   board[6][34] <= 0;
		   board[6][35] <= 0;
		   board[6][36] <= 0;
		   board[6][37] <= 0;
		   board[6][38] <= 0;
		   board[6][39] <= 0;
		   board[6][40] <= 0;
		   board[6][41] <= 0;
		   board[6][42] <= 0;
		   board[6][43] <= 0;
		   board[6][44] <= 0;
		   board[6][45] <= 0;
		   board[6][46] <= 0;
		   board[6][47] <= 0;
		   board[6][48] <= 0;
		   board[6][49] <= 0;
		   board[6][50] <= 0;
		   board[6][51] <= 0;
		   board[6][52] <= 0;
		   board[6][53] <= 0;
		   board[6][54] <= 0;
		   board[6][55] <= 0;
		   board[6][56] <= 0;
		   board[6][57] <= 0;
		   board[6][58] <= 0;
		   board[6][59] <= 0;
		   board[6][60] <= 0;
		   board[6][61] <= 0;
		   board[6][62] <= 0;
		   board[6][63] <= 0;
		   board[7][0] <= 0;
		   board[7][1] <= 0;
		   board[7][2] <= 0;
		   board[7][3] <= 0;
		   board[7][4] <= 0;
		   board[7][5] <= 0;
		   board[7][6] <= 0;
		   board[7][7] <= 0;
		   board[7][8] <= 0;
		   board[7][9] <= 0;
		   board[7][10] <= 0;
		   board[7][11] <= 0;
		   board[7][12] <= 0;
		   board[7][13] <= 0;
		   board[7][14] <= 0;
		   board[7][15] <= 0;
		   board[7][16] <= 0;
		   board[7][17] <= 0;
		   board[7][18] <= 0;
		   board[7][19] <= 0;
		   board[7][20] <= 0;
		   board[7][21] <= 0;
		   board[7][22] <= 0;
		   board[7][23] <= 0;
		   board[7][24] <= 0;
		   board[7][25] <= 0;
		   board[7][26] <= 0;
		   board[7][27] <= 0;
		   board[7][28] <= 0;
		   board[7][29] <= 0;
		   board[7][30] <= 0;
		   board[7][31] <= 0;
		   board[7][32] <= 0;
		   board[7][33] <= 0;
		   board[7][34] <= 0;
		   board[7][35] <= 0;
		   board[7][36] <= 0;
		   board[7][37] <= 0;
		   board[7][38] <= 0;
		   board[7][39] <= 0;
		   board[7][40] <= 0;
		   board[7][41] <= 0;
		   board[7][42] <= 0;
		   board[7][43] <= 0;
		   board[7][44] <= 0;
		   board[7][45] <= 0;
		   board[7][46] <= 0;
		   board[7][47] <= 0;
		   board[7][48] <= 0;
		   board[7][49] <= 0;
		   board[7][50] <= 0;
		   board[7][51] <= 0;
		   board[7][52] <= 0;
		   board[7][53] <= 0;
		   board[7][54] <= 0;
		   board[7][55] <= 0;
		   board[7][56] <= 0;
		   board[7][57] <= 0;
		   board[7][58] <= 0;
		   board[7][59] <= 0;
		   board[7][60] <= 0;
		   board[7][61] <= 0;
		   board[7][62] <= 0;
		   board[7][63] <= 0;
		   board[8][0] <= 0;
		   board[8][1] <= 0;
		   board[8][2] <= 0;
		   board[8][3] <= 0;
		   board[8][4] <= 0;
		   board[8][5] <= 0;
		   board[8][6] <= 0;
		   board[8][7] <= 0;
		   board[8][8] <= 0;
		   board[8][9] <= 0;
		   board[8][10] <= 0;
		   board[8][11] <= 0;
		   board[8][12] <= 0;
		   board[8][13] <= 0;
		   board[8][14] <= 0;
		   board[8][15] <= 0;
		   board[8][16] <= 0;
		   board[8][17] <= 0;
		   board[8][18] <= 0;
		   board[8][19] <= 0;
		   board[8][20] <= 0;
		   board[8][21] <= 0;
		   board[8][22] <= 0;
		   board[8][23] <= 0;
		   board[8][24] <= 0;
		   board[8][25] <= 0;
		   board[8][26] <= 0;
		   board[8][27] <= 0;
		   board[8][28] <= 0;
		   board[8][29] <= 0;
		   board[8][30] <= 0;
		   board[8][31] <= 0;
		   board[8][32] <= 0;
		   board[8][33] <= 0;
		   board[8][34] <= 0;
		   board[8][35] <= 0;
		   board[8][36] <= 0;
		   board[8][37] <= 0;
		   board[8][38] <= 0;
		   board[8][39] <= 0;
		   board[8][40] <= 0;
		   board[8][41] <= 0;
		   board[8][42] <= 0;
		   board[8][43] <= 0;
		   board[8][44] <= 0;
		   board[8][45] <= 0;
		   board[8][46] <= 0;
		   board[8][47] <= 0;
		   board[8][48] <= 0;
		   board[8][49] <= 0;
		   board[8][50] <= 0;
		   board[8][51] <= 0;
		   board[8][52] <= 0;
		   board[8][53] <= 0;
		   board[8][54] <= 0;
		   board[8][55] <= 0;
		   board[8][56] <= 0;
		   board[8][57] <= 0;
		   board[8][58] <= 0;
		   board[8][59] <= 0;
		   board[8][60] <= 0;
		   board[8][61] <= 0;
		   board[8][62] <= 0;
		   board[8][63] <= 0;
		   board[9][0] <= 0;
		   board[9][1] <= 0;
		   board[9][2] <= 0;
		   board[9][3] <= 0;
		   board[9][4] <= 0;
		   board[9][5] <= 0;
		   board[9][6] <= 0;
		   board[9][7] <= 0;
		   board[9][8] <= 0;
		   board[9][9] <= 0;
		   board[9][10] <= 0;
		   board[9][11] <= 0;
		   board[9][12] <= 0;
		   board[9][13] <= 0;
		   board[9][14] <= 0;
		   board[9][15] <= 0;
		   board[9][16] <= 0;
		   board[9][17] <= 0;
		   board[9][18] <= 0;
		   board[9][19] <= 0;
		   board[9][20] <= 0;
		   board[9][21] <= 0;
		   board[9][22] <= 0;
		   board[9][23] <= 0;
		   board[9][24] <= 0;
		   board[9][25] <= 0;
		   board[9][26] <= 0;
		   board[9][27] <= 0;
		   board[9][28] <= 0;
		   board[9][29] <= 0;
		   board[9][30] <= 0;
		   board[9][31] <= 1;
		   board[9][32] <= 0;
		   board[9][33] <= 0;
		   board[9][34] <= 0;
		   board[9][35] <= 0;
		   board[9][36] <= 0;
		   board[9][37] <= 0;
		   board[9][38] <= 0;
		   board[9][39] <= 0;
		   board[9][40] <= 0;
		   board[9][41] <= 0;
		   board[9][42] <= 0;
		   board[9][43] <= 0;
		   board[9][44] <= 0;
		   board[9][45] <= 0;
		   board[9][46] <= 0;
		   board[9][47] <= 0;
		   board[9][48] <= 0;
		   board[9][49] <= 0;
		   board[9][50] <= 0;
		   board[9][51] <= 0;
		   board[9][52] <= 0;
		   board[9][53] <= 0;
		   board[9][54] <= 0;
		   board[9][55] <= 0;
		   board[9][56] <= 0;
		   board[9][57] <= 0;
		   board[9][58] <= 0;
		   board[9][59] <= 0;
		   board[9][60] <= 0;
		   board[9][61] <= 0;
		   board[9][62] <= 0;
		   board[9][63] <= 0;
		   board[10][0] <= 0;
		   board[10][1] <= 0;
		   board[10][2] <= 0;
		   board[10][3] <= 0;
		   board[10][4] <= 0;
		   board[10][5] <= 0;
		   board[10][6] <= 0;
		   board[10][7] <= 0;
		   board[10][8] <= 0;
		   board[10][9] <= 0;
		   board[10][10] <= 0;
		   board[10][11] <= 0;
		   board[10][12] <= 0;
		   board[10][13] <= 0;
		   board[10][14] <= 0;
		   board[10][15] <= 0;
		   board[10][16] <= 0;
		   board[10][17] <= 0;
		   board[10][18] <= 0;
		   board[10][19] <= 0;
		   board[10][20] <= 0;
		   board[10][21] <= 0;
		   board[10][22] <= 0;
		   board[10][23] <= 0;
		   board[10][24] <= 0;
		   board[10][25] <= 0;
		   board[10][26] <= 0;
		   board[10][27] <= 0;
		   board[10][28] <= 0;
		   board[10][29] <= 1;
		   board[10][30] <= 0;
		   board[10][31] <= 1;
		   board[10][32] <= 0;
		   board[10][33] <= 0;
		   board[10][34] <= 0;
		   board[10][35] <= 0;
		   board[10][36] <= 0;
		   board[10][37] <= 0;
		   board[10][38] <= 0;
		   board[10][39] <= 0;
		   board[10][40] <= 0;
		   board[10][41] <= 0;
		   board[10][42] <= 0;
		   board[10][43] <= 0;
		   board[10][44] <= 0;
		   board[10][45] <= 0;
		   board[10][46] <= 0;
		   board[10][47] <= 0;
		   board[10][48] <= 0;
		   board[10][49] <= 0;
		   board[10][50] <= 0;
		   board[10][51] <= 0;
		   board[10][52] <= 0;
		   board[10][53] <= 0;
		   board[10][54] <= 0;
		   board[10][55] <= 0;
		   board[10][56] <= 0;
		   board[10][57] <= 0;
		   board[10][58] <= 0;
		   board[10][59] <= 0;
		   board[10][60] <= 0;
		   board[10][61] <= 0;
		   board[10][62] <= 0;
		   board[10][63] <= 0;
		   board[11][0] <= 0;
		   board[11][1] <= 0;
		   board[11][2] <= 0;
		   board[11][3] <= 0;
		   board[11][4] <= 0;
		   board[11][5] <= 0;
		   board[11][6] <= 0;
		   board[11][7] <= 0;
		   board[11][8] <= 0;
		   board[11][9] <= 0;
		   board[11][10] <= 0;
		   board[11][11] <= 0;
		   board[11][12] <= 0;
		   board[11][13] <= 0;
		   board[11][14] <= 0;
		   board[11][15] <= 0;
		   board[11][16] <= 0;
		   board[11][17] <= 0;
		   board[11][18] <= 0;
		   board[11][19] <= 1;
		   board[11][20] <= 1;
		   board[11][21] <= 0;
		   board[11][22] <= 0;
		   board[11][23] <= 0;
		   board[11][24] <= 0;
		   board[11][25] <= 0;
		   board[11][26] <= 0;
		   board[11][27] <= 1;
		   board[11][28] <= 1;
		   board[11][29] <= 0;
		   board[11][30] <= 0;
		   board[11][31] <= 0;
		   board[11][32] <= 0;
		   board[11][33] <= 0;
		   board[11][34] <= 0;
		   board[11][35] <= 0;
		   board[11][36] <= 0;
		   board[11][37] <= 0;
		   board[11][38] <= 0;
		   board[11][39] <= 0;
		   board[11][40] <= 0;
		   board[11][41] <= 1;
		   board[11][42] <= 1;
		   board[11][43] <= 0;
		   board[11][44] <= 0;
		   board[11][45] <= 0;
		   board[11][46] <= 0;
		   board[11][47] <= 0;
		   board[11][48] <= 0;
		   board[11][49] <= 0;
		   board[11][50] <= 0;
		   board[11][51] <= 0;
		   board[11][52] <= 0;
		   board[11][53] <= 0;
		   board[11][54] <= 0;
		   board[11][55] <= 0;
		   board[11][56] <= 0;
		   board[11][57] <= 0;
		   board[11][58] <= 0;
		   board[11][59] <= 0;
		   board[11][60] <= 0;
		   board[11][61] <= 0;
		   board[11][62] <= 0;
		   board[11][63] <= 0;
		   board[12][0] <= 0;
		   board[12][1] <= 0;
		   board[12][2] <= 0;
		   board[12][3] <= 0;
		   board[12][4] <= 0;
		   board[12][5] <= 0;
		   board[12][6] <= 0;
		   board[12][7] <= 0;
		   board[12][8] <= 0;
		   board[12][9] <= 0;
		   board[12][10] <= 0;
		   board[12][11] <= 0;
		   board[12][12] <= 0;
		   board[12][13] <= 0;
		   board[12][14] <= 0;
		   board[12][15] <= 0;
		   board[12][16] <= 0;
		   board[12][17] <= 0;
		   board[12][18] <= 1;
		   board[12][19] <= 0;
		   board[12][20] <= 0;
		   board[12][21] <= 0;
		   board[12][22] <= 1;
		   board[12][23] <= 0;
		   board[12][24] <= 0;
		   board[12][25] <= 0;
		   board[12][26] <= 0;
		   board[12][27] <= 1;
		   board[12][28] <= 1;
		   board[12][29] <= 0;
		   board[12][30] <= 0;
		   board[12][31] <= 0;
		   board[12][32] <= 0;
		   board[12][33] <= 0;
		   board[12][34] <= 0;
		   board[12][35] <= 0;
		   board[12][36] <= 0;
		   board[12][37] <= 0;
		   board[12][38] <= 0;
		   board[12][39] <= 0;
		   board[12][40] <= 0;
		   board[12][41] <= 1;
		   board[12][42] <= 1;
		   board[12][43] <= 0;
		   board[12][44] <= 0;
		   board[12][45] <= 0;
		   board[12][46] <= 0;
		   board[12][47] <= 0;
		   board[12][48] <= 0;
		   board[12][49] <= 0;
		   board[12][50] <= 0;
		   board[12][51] <= 0;
		   board[12][52] <= 0;
		   board[12][53] <= 0;
		   board[12][54] <= 0;
		   board[12][55] <= 0;
		   board[12][56] <= 0;
		   board[12][57] <= 0;
		   board[12][58] <= 0;
		   board[12][59] <= 0;
		   board[12][60] <= 0;
		   board[12][61] <= 0;
		   board[12][62] <= 0;
		   board[12][63] <= 0;
		   board[13][0] <= 0;
		   board[13][1] <= 0;
		   board[13][2] <= 0;
		   board[13][3] <= 0;
		   board[13][4] <= 0;
		   board[13][5] <= 0;
		   board[13][6] <= 0;
		   board[13][7] <= 1;
		   board[13][8] <= 1;
		   board[13][9] <= 0;
		   board[13][10] <= 0;
		   board[13][11] <= 0;
		   board[13][12] <= 0;
		   board[13][13] <= 0;
		   board[13][14] <= 0;
		   board[13][15] <= 0;
		   board[13][16] <= 0;
		   board[13][17] <= 1;
		   board[13][18] <= 0;
		   board[13][19] <= 0;
		   board[13][20] <= 0;
		   board[13][21] <= 0;
		   board[13][22] <= 0;
		   board[13][23] <= 1;
		   board[13][24] <= 0;
		   board[13][25] <= 0;
		   board[13][26] <= 0;
		   board[13][27] <= 1;
		   board[13][28] <= 1;
		   board[13][29] <= 0;
		   board[13][30] <= 0;
		   board[13][31] <= 0;
		   board[13][32] <= 0;
		   board[13][33] <= 0;
		   board[13][34] <= 0;
		   board[13][35] <= 0;
		   board[13][36] <= 0;
		   board[13][37] <= 0;
		   board[13][38] <= 0;
		   board[13][39] <= 0;
		   board[13][40] <= 0;
		   board[13][41] <= 0;
		   board[13][42] <= 0;
		   board[13][43] <= 0;
		   board[13][44] <= 0;
		   board[13][45] <= 0;
		   board[13][46] <= 0;
		   board[13][47] <= 0;
		   board[13][48] <= 0;
		   board[13][49] <= 0;
		   board[13][50] <= 0;
		   board[13][51] <= 0;
		   board[13][52] <= 0;
		   board[13][53] <= 0;
		   board[13][54] <= 0;
		   board[13][55] <= 0;
		   board[13][56] <= 0;
		   board[13][57] <= 0;
		   board[13][58] <= 0;
		   board[13][59] <= 0;
		   board[13][60] <= 0;
		   board[13][61] <= 0;
		   board[13][62] <= 0;
		   board[13][63] <= 0;
		   board[14][0] <= 0;
		   board[14][1] <= 0;
		   board[14][2] <= 0;
		   board[14][3] <= 0;
		   board[14][4] <= 0;
		   board[14][5] <= 0;
		   board[14][6] <= 0;
		   board[14][7] <= 1;
		   board[14][8] <= 1;
		   board[14][9] <= 0;
		   board[14][10] <= 0;
		   board[14][11] <= 0;
		   board[14][12] <= 0;
		   board[14][13] <= 0;
		   board[14][14] <= 0;
		   board[14][15] <= 0;
		   board[14][16] <= 0;
		   board[14][17] <= 1;
		   board[14][18] <= 0;
		   board[14][19] <= 0;
		   board[14][20] <= 0;
		   board[14][21] <= 1;
		   board[14][22] <= 0;
		   board[14][23] <= 1;
		   board[14][24] <= 1;
		   board[14][25] <= 0;
		   board[14][26] <= 0;
		   board[14][27] <= 0;
		   board[14][28] <= 0;
		   board[14][29] <= 1;
		   board[14][30] <= 0;
		   board[14][31] <= 1;
		   board[14][32] <= 0;
		   board[14][33] <= 0;
		   board[14][34] <= 0;
		   board[14][35] <= 0;
		   board[14][36] <= 0;
		   board[14][37] <= 0;
		   board[14][38] <= 0;
		   board[14][39] <= 0;
		   board[14][40] <= 0;
		   board[14][41] <= 0;
		   board[14][42] <= 0;
		   board[14][43] <= 0;
		   board[14][44] <= 0;
		   board[14][45] <= 0;
		   board[14][46] <= 0;
		   board[14][47] <= 0;
		   board[14][48] <= 0;
		   board[14][49] <= 0;
		   board[14][50] <= 0;
		   board[14][51] <= 0;
		   board[14][52] <= 0;
		   board[14][53] <= 0;
		   board[14][54] <= 0;
		   board[14][55] <= 0;
		   board[14][56] <= 0;
		   board[14][57] <= 0;
		   board[14][58] <= 0;
		   board[14][59] <= 0;
		   board[14][60] <= 0;
		   board[14][61] <= 0;
		   board[14][62] <= 0;
		   board[14][63] <= 0;
		   board[15][0] <= 0;
		   board[15][1] <= 0;
		   board[15][2] <= 0;
		   board[15][3] <= 0;
		   board[15][4] <= 0;
		   board[15][5] <= 0;
		   board[15][6] <= 0;
		   board[15][7] <= 0;
		   board[15][8] <= 0;
		   board[15][9] <= 0;
		   board[15][10] <= 0;
		   board[15][11] <= 0;
		   board[15][12] <= 0;
		   board[15][13] <= 0;
		   board[15][14] <= 0;
		   board[15][15] <= 0;
		   board[15][16] <= 0;
		   board[15][17] <= 1;
		   board[15][18] <= 0;
		   board[15][19] <= 0;
		   board[15][20] <= 0;
		   board[15][21] <= 0;
		   board[15][22] <= 0;
		   board[15][23] <= 1;
		   board[15][24] <= 0;
		   board[15][25] <= 0;
		   board[15][26] <= 0;
		   board[15][27] <= 0;
		   board[15][28] <= 0;
		   board[15][29] <= 0;
		   board[15][30] <= 0;
		   board[15][31] <= 1;
		   board[15][32] <= 0;
		   board[15][33] <= 0;
		   board[15][34] <= 0;
		   board[15][35] <= 0;
		   board[15][36] <= 0;
		   board[15][37] <= 0;
		   board[15][38] <= 0;
		   board[15][39] <= 0;
		   board[15][40] <= 0;
		   board[15][41] <= 0;
		   board[15][42] <= 0;
		   board[15][43] <= 0;
		   board[15][44] <= 0;
		   board[15][45] <= 0;
		   board[15][46] <= 0;
		   board[15][47] <= 0;
		   board[15][48] <= 0;
		   board[15][49] <= 0;
		   board[15][50] <= 0;
		   board[15][51] <= 0;
		   board[15][52] <= 0;
		   board[15][53] <= 0;
		   board[15][54] <= 0;
		   board[15][55] <= 0;
		   board[15][56] <= 0;
		   board[15][57] <= 0;
		   board[15][58] <= 0;
		   board[15][59] <= 0;
		   board[15][60] <= 0;
		   board[15][61] <= 0;
		   board[15][62] <= 0;
		   board[15][63] <= 0;
		   board[16][0] <= 0;
		   board[16][1] <= 0;
		   board[16][2] <= 0;
		   board[16][3] <= 0;
		   board[16][4] <= 0;
		   board[16][5] <= 0;
		   board[16][6] <= 0;
		   board[16][7] <= 0;
		   board[16][8] <= 0;
		   board[16][9] <= 0;
		   board[16][10] <= 0;
		   board[16][11] <= 0;
		   board[16][12] <= 0;
		   board[16][13] <= 0;
		   board[16][14] <= 0;
		   board[16][15] <= 0;
		   board[16][16] <= 0;
		   board[16][17] <= 0;
		   board[16][18] <= 1;
		   board[16][19] <= 0;
		   board[16][20] <= 0;
		   board[16][21] <= 0;
		   board[16][22] <= 1;
		   board[16][23] <= 0;
		   board[16][24] <= 0;
		   board[16][25] <= 0;
		   board[16][26] <= 0;
		   board[16][27] <= 0;
		   board[16][28] <= 0;
		   board[16][29] <= 0;
		   board[16][30] <= 0;
		   board[16][31] <= 0;
		   board[16][32] <= 0;
		   board[16][33] <= 0;
		   board[16][34] <= 0;
		   board[16][35] <= 0;
		   board[16][36] <= 0;
		   board[16][37] <= 0;
		   board[16][38] <= 0;
		   board[16][39] <= 0;
		   board[16][40] <= 0;
		   board[16][41] <= 0;
		   board[16][42] <= 0;
		   board[16][43] <= 0;
		   board[16][44] <= 0;
		   board[16][45] <= 0;
		   board[16][46] <= 0;
		   board[16][47] <= 0;
		   board[16][48] <= 0;
		   board[16][49] <= 0;
		   board[16][50] <= 0;
		   board[16][51] <= 0;
		   board[16][52] <= 0;
		   board[16][53] <= 0;
		   board[16][54] <= 0;
		   board[16][55] <= 0;
		   board[16][56] <= 0;
		   board[16][57] <= 0;
		   board[16][58] <= 0;
		   board[16][59] <= 0;
		   board[16][60] <= 0;
		   board[16][61] <= 0;
		   board[16][62] <= 0;
		   board[16][63] <= 0;
		   board[17][0] <= 0;
		   board[17][1] <= 0;
		   board[17][2] <= 0;
		   board[17][3] <= 0;
		   board[17][4] <= 0;
		   board[17][5] <= 0;
		   board[17][6] <= 0;
		   board[17][7] <= 0;
		   board[17][8] <= 0;
		   board[17][9] <= 0;
		   board[17][10] <= 0;
		   board[17][11] <= 0;
		   board[17][12] <= 0;
		   board[17][13] <= 0;
		   board[17][14] <= 0;
		   board[17][15] <= 0;
		   board[17][16] <= 0;
		   board[17][17] <= 0;
		   board[17][18] <= 0;
		   board[17][19] <= 1;
		   board[17][20] <= 1;
		   board[17][21] <= 0;
		   board[17][22] <= 0;
		   board[17][23] <= 0;
		   board[17][24] <= 0;
		   board[17][25] <= 0;
		   board[17][26] <= 0;
		   board[17][27] <= 0;
		   board[17][28] <= 0;
		   board[17][29] <= 0;
		   board[17][30] <= 0;
		   board[17][31] <= 0;
		   board[17][32] <= 0;
		   board[17][33] <= 0;
		   board[17][34] <= 0;
		   board[17][35] <= 0;
		   board[17][36] <= 0;
		   board[17][37] <= 0;
		   board[17][38] <= 0;
		   board[17][39] <= 0;
		   board[17][40] <= 0;
		   board[17][41] <= 0;
		   board[17][42] <= 0;
		   board[17][43] <= 0;
		   board[17][44] <= 0;
		   board[17][45] <= 0;
		   board[17][46] <= 0;
		   board[17][47] <= 0;
		   board[17][48] <= 0;
		   board[17][49] <= 0;
		   board[17][50] <= 0;
		   board[17][51] <= 0;
		   board[17][52] <= 0;
		   board[17][53] <= 0;
		   board[17][54] <= 0;
		   board[17][55] <= 0;
		   board[17][56] <= 0;
		   board[17][57] <= 0;
		   board[17][58] <= 0;
		   board[17][59] <= 0;
		   board[17][60] <= 0;
		   board[17][61] <= 0;
		   board[17][62] <= 0;
		   board[17][63] <= 0;
		   board[18][0] <= 0;
		   board[18][1] <= 0;
		   board[18][2] <= 0;
		   board[18][3] <= 0;
		   board[18][4] <= 0;
		   board[18][5] <= 0;
		   board[18][6] <= 0;
		   board[18][7] <= 0;
		   board[18][8] <= 0;
		   board[18][9] <= 0;
		   board[18][10] <= 0;
		   board[18][11] <= 0;
		   board[18][12] <= 0;
		   board[18][13] <= 0;
		   board[18][14] <= 0;
		   board[18][15] <= 0;
		   board[18][16] <= 0;
		   board[18][17] <= 0;
		   board[18][18] <= 0;
		   board[18][19] <= 0;
		   board[18][20] <= 0;
		   board[18][21] <= 0;
		   board[18][22] <= 0;
		   board[18][23] <= 0;
		   board[18][24] <= 0;
		   board[18][25] <= 0;
		   board[18][26] <= 0;
		   board[18][27] <= 0;
		   board[18][28] <= 0;
		   board[18][29] <= 0;
		   board[18][30] <= 0;
		   board[18][31] <= 0;
		   board[18][32] <= 0;
		   board[18][33] <= 0;
		   board[18][34] <= 0;
		   board[18][35] <= 0;
		   board[18][36] <= 0;
		   board[18][37] <= 0;
		   board[18][38] <= 0;
		   board[18][39] <= 0;
		   board[18][40] <= 0;
		   board[18][41] <= 0;
		   board[18][42] <= 0;
		   board[18][43] <= 0;
		   board[18][44] <= 0;
		   board[18][45] <= 0;
		   board[18][46] <= 0;
		   board[18][47] <= 0;
		   board[18][48] <= 0;
		   board[18][49] <= 0;
		   board[18][50] <= 0;
		   board[18][51] <= 0;
		   board[18][52] <= 0;
		   board[18][53] <= 0;
		   board[18][54] <= 0;
		   board[18][55] <= 0;
		   board[18][56] <= 0;
		   board[18][57] <= 0;
		   board[18][58] <= 0;
		   board[18][59] <= 0;
		   board[18][60] <= 0;
		   board[18][61] <= 0;
		   board[18][62] <= 0;
		   board[18][63] <= 0;
		   board[19][0] <= 0;
		   board[19][1] <= 0;
		   board[19][2] <= 0;
		   board[19][3] <= 0;
		   board[19][4] <= 0;
		   board[19][5] <= 0;
		   board[19][6] <= 0;
		   board[19][7] <= 0;
		   board[19][8] <= 0;
		   board[19][9] <= 0;
		   board[19][10] <= 0;
		   board[19][11] <= 0;
		   board[19][12] <= 0;
		   board[19][13] <= 0;
		   board[19][14] <= 0;
		   board[19][15] <= 0;
		   board[19][16] <= 0;
		   board[19][17] <= 0;
		   board[19][18] <= 0;
		   board[19][19] <= 0;
		   board[19][20] <= 0;
		   board[19][21] <= 0;
		   board[19][22] <= 0;
		   board[19][23] <= 0;
		   board[19][24] <= 0;
		   board[19][25] <= 0;
		   board[19][26] <= 0;
		   board[19][27] <= 0;
		   board[19][28] <= 0;
		   board[19][29] <= 0;
		   board[19][30] <= 0;
		   board[19][31] <= 0;
		   board[19][32] <= 0;
		   board[19][33] <= 0;
		   board[19][34] <= 0;
		   board[19][35] <= 0;
		   board[19][36] <= 0;
		   board[19][37] <= 0;
		   board[19][38] <= 0;
		   board[19][39] <= 0;
		   board[19][40] <= 0;
		   board[19][41] <= 0;
		   board[19][42] <= 0;
		   board[19][43] <= 0;
		   board[19][44] <= 0;
		   board[19][45] <= 0;
		   board[19][46] <= 0;
		   board[19][47] <= 0;
		   board[19][48] <= 0;
		   board[19][49] <= 0;
		   board[19][50] <= 0;
		   board[19][51] <= 0;
		   board[19][52] <= 0;
		   board[19][53] <= 0;
		   board[19][54] <= 0;
		   board[19][55] <= 0;
		   board[19][56] <= 0;
		   board[19][57] <= 0;
		   board[19][58] <= 0;
		   board[19][59] <= 0;
		   board[19][60] <= 0;
		   board[19][61] <= 0;
		   board[19][62] <= 0;
		   board[19][63] <= 0;
		   board[20][0] <= 0;
		   board[20][1] <= 0;
		   board[20][2] <= 0;
		   board[20][3] <= 0;
		   board[20][4] <= 0;
		   board[20][5] <= 0;
		   board[20][6] <= 0;
		   board[20][7] <= 0;
		   board[20][8] <= 0;
		   board[20][9] <= 0;
		   board[20][10] <= 0;
		   board[20][11] <= 0;
		   board[20][12] <= 0;
		   board[20][13] <= 0;
		   board[20][14] <= 0;
		   board[20][15] <= 0;
		   board[20][16] <= 0;
		   board[20][17] <= 0;
		   board[20][18] <= 0;
		   board[20][19] <= 0;
		   board[20][20] <= 0;
		   board[20][21] <= 0;
		   board[20][22] <= 0;
		   board[20][23] <= 0;
		   board[20][24] <= 0;
		   board[20][25] <= 0;
		   board[20][26] <= 0;
		   board[20][27] <= 0;
		   board[20][28] <= 0;
		   board[20][29] <= 0;
		   board[20][30] <= 0;
		   board[20][31] <= 0;
		   board[20][32] <= 0;
		   board[20][33] <= 0;
		   board[20][34] <= 0;
		   board[20][35] <= 0;
		   board[20][36] <= 0;
		   board[20][37] <= 0;
		   board[20][38] <= 0;
		   board[20][39] <= 0;
		   board[20][40] <= 0;
		   board[20][41] <= 0;
		   board[20][42] <= 0;
		   board[20][43] <= 0;
		   board[20][44] <= 0;
		   board[20][45] <= 0;
		   board[20][46] <= 0;
		   board[20][47] <= 0;
		   board[20][48] <= 0;
		   board[20][49] <= 0;
		   board[20][50] <= 0;
		   board[20][51] <= 0;
		   board[20][52] <= 0;
		   board[20][53] <= 0;
		   board[20][54] <= 0;
		   board[20][55] <= 0;
		   board[20][56] <= 0;
		   board[20][57] <= 0;
		   board[20][58] <= 0;
		   board[20][59] <= 0;
		   board[20][60] <= 0;
		   board[20][61] <= 0;
		   board[20][62] <= 0;
		   board[20][63] <= 0;
		   board[21][0] <= 0;
		   board[21][1] <= 0;
		   board[21][2] <= 0;
		   board[21][3] <= 0;
		   board[21][4] <= 0;
		   board[21][5] <= 0;
		   board[21][6] <= 0;
		   board[21][7] <= 0;
		   board[21][8] <= 0;
		   board[21][9] <= 0;
		   board[21][10] <= 0;
		   board[21][11] <= 0;
		   board[21][12] <= 0;
		   board[21][13] <= 0;
		   board[21][14] <= 0;
		   board[21][15] <= 0;
		   board[21][16] <= 0;
		   board[21][17] <= 0;
		   board[21][18] <= 0;
		   board[21][19] <= 0;
		   board[21][20] <= 0;
		   board[21][21] <= 0;
		   board[21][22] <= 0;
		   board[21][23] <= 0;
		   board[21][24] <= 0;
		   board[21][25] <= 0;
		   board[21][26] <= 0;
		   board[21][27] <= 0;
		   board[21][28] <= 0;
		   board[21][29] <= 0;
		   board[21][30] <= 0;
		   board[21][31] <= 0;
		   board[21][32] <= 0;
		   board[21][33] <= 0;
		   board[21][34] <= 0;
		   board[21][35] <= 0;
		   board[21][36] <= 0;
		   board[21][37] <= 0;
		   board[21][38] <= 0;
		   board[21][39] <= 0;
		   board[21][40] <= 0;
		   board[21][41] <= 0;
		   board[21][42] <= 0;
		   board[21][43] <= 0;
		   board[21][44] <= 0;
		   board[21][45] <= 0;
		   board[21][46] <= 0;
		   board[21][47] <= 0;
		   board[21][48] <= 0;
		   board[21][49] <= 0;
		   board[21][50] <= 0;
		   board[21][51] <= 0;
		   board[21][52] <= 0;
		   board[21][53] <= 0;
		   board[21][54] <= 0;
		   board[21][55] <= 0;
		   board[21][56] <= 0;
		   board[21][57] <= 0;
		   board[21][58] <= 0;
		   board[21][59] <= 0;
		   board[21][60] <= 0;
		   board[21][61] <= 0;
		   board[21][62] <= 0;
		   board[21][63] <= 0;
		   board[22][0] <= 0;
		   board[22][1] <= 0;
		   board[22][2] <= 0;
		   board[22][3] <= 0;
		   board[22][4] <= 0;
		   board[22][5] <= 0;
		   board[22][6] <= 0;
		   board[22][7] <= 0;
		   board[22][8] <= 0;
		   board[22][9] <= 0;
		   board[22][10] <= 0;
		   board[22][11] <= 0;
		   board[22][12] <= 0;
		   board[22][13] <= 0;
		   board[22][14] <= 0;
		   board[22][15] <= 0;
		   board[22][16] <= 0;
		   board[22][17] <= 0;
		   board[22][18] <= 0;
		   board[22][19] <= 0;
		   board[22][20] <= 0;
		   board[22][21] <= 0;
		   board[22][22] <= 0;
		   board[22][23] <= 0;
		   board[22][24] <= 0;
		   board[22][25] <= 0;
		   board[22][26] <= 0;
		   board[22][27] <= 0;
		   board[22][28] <= 0;
		   board[22][29] <= 0;
		   board[22][30] <= 0;
		   board[22][31] <= 0;
		   board[22][32] <= 0;
		   board[22][33] <= 0;
		   board[22][34] <= 0;
		   board[22][35] <= 0;
		   board[22][36] <= 0;
		   board[22][37] <= 0;
		   board[22][38] <= 0;
		   board[22][39] <= 0;
		   board[22][40] <= 0;
		   board[22][41] <= 0;
		   board[22][42] <= 0;
		   board[22][43] <= 0;
		   board[22][44] <= 0;
		   board[22][45] <= 0;
		   board[22][46] <= 0;
		   board[22][47] <= 0;
		   board[22][48] <= 0;
		   board[22][49] <= 0;
		   board[22][50] <= 0;
		   board[22][51] <= 0;
		   board[22][52] <= 0;
		   board[22][53] <= 0;
		   board[22][54] <= 0;
		   board[22][55] <= 0;
		   board[22][56] <= 0;
		   board[22][57] <= 0;
		   board[22][58] <= 0;
		   board[22][59] <= 0;
		   board[22][60] <= 0;
		   board[22][61] <= 0;
		   board[22][62] <= 0;
		   board[22][63] <= 0;
		   board[23][0] <= 0;
		   board[23][1] <= 0;
		   board[23][2] <= 0;
		   board[23][3] <= 0;
		   board[23][4] <= 0;
		   board[23][5] <= 0;
		   board[23][6] <= 0;
		   board[23][7] <= 0;
		   board[23][8] <= 0;
		   board[23][9] <= 0;
		   board[23][10] <= 0;
		   board[23][11] <= 0;
		   board[23][12] <= 0;
		   board[23][13] <= 0;
		   board[23][14] <= 0;
		   board[23][15] <= 0;
		   board[23][16] <= 0;
		   board[23][17] <= 0;
		   board[23][18] <= 0;
		   board[23][19] <= 0;
		   board[23][20] <= 0;
		   board[23][21] <= 0;
		   board[23][22] <= 0;
		   board[23][23] <= 0;
		   board[23][24] <= 0;
		   board[23][25] <= 0;
		   board[23][26] <= 0;
		   board[23][27] <= 0;
		   board[23][28] <= 0;
		   board[23][29] <= 0;
		   board[23][30] <= 0;
		   board[23][31] <= 0;
		   board[23][32] <= 0;
		   board[23][33] <= 0;
		   board[23][34] <= 0;
		   board[23][35] <= 0;
		   board[23][36] <= 0;
		   board[23][37] <= 0;
		   board[23][38] <= 0;
		   board[23][39] <= 0;
		   board[23][40] <= 0;
		   board[23][41] <= 0;
		   board[23][42] <= 0;
		   board[23][43] <= 0;
		   board[23][44] <= 0;
		   board[23][45] <= 0;
		   board[23][46] <= 0;
		   board[23][47] <= 0;
		   board[23][48] <= 0;
		   board[23][49] <= 0;
		   board[23][50] <= 0;
		   board[23][51] <= 0;
		   board[23][52] <= 0;
		   board[23][53] <= 0;
		   board[23][54] <= 0;
		   board[23][55] <= 0;
		   board[23][56] <= 0;
		   board[23][57] <= 0;
		   board[23][58] <= 0;
		   board[23][59] <= 0;
		   board[23][60] <= 0;
		   board[23][61] <= 0;
		   board[23][62] <= 0;
		   board[23][63] <= 0;
		   board[24][0] <= 0;
		   board[24][1] <= 0;
		   board[24][2] <= 0;
		   board[24][3] <= 0;
		   board[24][4] <= 0;
		   board[24][5] <= 0;
		   board[24][6] <= 0;
		   board[24][7] <= 0;
		   board[24][8] <= 0;
		   board[24][9] <= 0;
		   board[24][10] <= 0;
		   board[24][11] <= 0;
		   board[24][12] <= 0;
		   board[24][13] <= 0;
		   board[24][14] <= 0;
		   board[24][15] <= 0;
		   board[24][16] <= 0;
		   board[24][17] <= 0;
		   board[24][18] <= 0;
		   board[24][19] <= 0;
		   board[24][20] <= 0;
		   board[24][21] <= 0;
		   board[24][22] <= 0;
		   board[24][23] <= 0;
		   board[24][24] <= 0;
		   board[24][25] <= 0;
		   board[24][26] <= 0;
		   board[24][27] <= 0;
		   board[24][28] <= 0;
		   board[24][29] <= 0;
		   board[24][30] <= 0;
		   board[24][31] <= 0;
		   board[24][32] <= 0;
		   board[24][33] <= 0;
		   board[24][34] <= 0;
		   board[24][35] <= 0;
		   board[24][36] <= 0;
		   board[24][37] <= 0;
		   board[24][38] <= 0;
		   board[24][39] <= 0;
		   board[24][40] <= 0;
		   board[24][41] <= 0;
		   board[24][42] <= 0;
		   board[24][43] <= 0;
		   board[24][44] <= 0;
		   board[24][45] <= 0;
		   board[24][46] <= 0;
		   board[24][47] <= 0;
		   board[24][48] <= 0;
		   board[24][49] <= 0;
		   board[24][50] <= 0;
		   board[24][51] <= 0;
		   board[24][52] <= 0;
		   board[24][53] <= 0;
		   board[24][54] <= 0;
		   board[24][55] <= 0;
		   board[24][56] <= 0;
		   board[24][57] <= 0;
		   board[24][58] <= 0;
		   board[24][59] <= 0;
		   board[24][60] <= 0;
		   board[24][61] <= 0;
		   board[24][62] <= 0;
		   board[24][63] <= 0;
		   board[25][0] <= 0;
		   board[25][1] <= 0;
		   board[25][2] <= 0;
		   board[25][3] <= 0;
		   board[25][4] <= 0;
		   board[25][5] <= 0;
		   board[25][6] <= 0;
		   board[25][7] <= 0;
		   board[25][8] <= 0;
		   board[25][9] <= 0;
		   board[25][10] <= 0;
		   board[25][11] <= 0;
		   board[25][12] <= 0;
		   board[25][13] <= 0;
		   board[25][14] <= 0;
		   board[25][15] <= 0;
		   board[25][16] <= 0;
		   board[25][17] <= 0;
		   board[25][18] <= 0;
		   board[25][19] <= 0;
		   board[25][20] <= 0;
		   board[25][21] <= 0;
		   board[25][22] <= 0;
		   board[25][23] <= 0;
		   board[25][24] <= 0;
		   board[25][25] <= 0;
		   board[25][26] <= 0;
		   board[25][27] <= 0;
		   board[25][28] <= 0;
		   board[25][29] <= 0;
		   board[25][30] <= 0;
		   board[25][31] <= 0;
		   board[25][32] <= 0;
		   board[25][33] <= 0;
		   board[25][34] <= 0;
		   board[25][35] <= 0;
		   board[25][36] <= 0;
		   board[25][37] <= 0;
		   board[25][38] <= 0;
		   board[25][39] <= 0;
		   board[25][40] <= 0;
		   board[25][41] <= 0;
		   board[25][42] <= 0;
		   board[25][43] <= 0;
		   board[25][44] <= 0;
		   board[25][45] <= 0;
		   board[25][46] <= 0;
		   board[25][47] <= 0;
		   board[25][48] <= 0;
		   board[25][49] <= 0;
		   board[25][50] <= 0;
		   board[25][51] <= 0;
		   board[25][52] <= 0;
		   board[25][53] <= 0;
		   board[25][54] <= 0;
		   board[25][55] <= 0;
		   board[25][56] <= 0;
		   board[25][57] <= 0;
		   board[25][58] <= 0;
		   board[25][59] <= 0;
		   board[25][60] <= 0;
		   board[25][61] <= 0;
		   board[25][62] <= 0;
		   board[25][63] <= 0;
		   board[26][0] <= 0;
		   board[26][1] <= 0;
		   board[26][2] <= 0;
		   board[26][3] <= 0;
		   board[26][4] <= 0;
		   board[26][5] <= 0;
		   board[26][6] <= 0;
		   board[26][7] <= 0;
		   board[26][8] <= 0;
		   board[26][9] <= 0;
		   board[26][10] <= 0;
		   board[26][11] <= 0;
		   board[26][12] <= 0;
		   board[26][13] <= 0;
		   board[26][14] <= 0;
		   board[26][15] <= 0;
		   board[26][16] <= 0;
		   board[26][17] <= 0;
		   board[26][18] <= 0;
		   board[26][19] <= 0;
		   board[26][20] <= 0;
		   board[26][21] <= 0;
		   board[26][22] <= 0;
		   board[26][23] <= 0;
		   board[26][24] <= 0;
		   board[26][25] <= 0;
		   board[26][26] <= 0;
		   board[26][27] <= 0;
		   board[26][28] <= 0;
		   board[26][29] <= 0;
		   board[26][30] <= 0;
		   board[26][31] <= 0;
		   board[26][32] <= 0;
		   board[26][33] <= 0;
		   board[26][34] <= 0;
		   board[26][35] <= 0;
		   board[26][36] <= 0;
		   board[26][37] <= 0;
		   board[26][38] <= 0;
		   board[26][39] <= 0;
		   board[26][40] <= 0;
		   board[26][41] <= 0;
		   board[26][42] <= 0;
		   board[26][43] <= 0;
		   board[26][44] <= 0;
		   board[26][45] <= 0;
		   board[26][46] <= 0;
		   board[26][47] <= 0;
		   board[26][48] <= 0;
		   board[26][49] <= 0;
		   board[26][50] <= 0;
		   board[26][51] <= 0;
		   board[26][52] <= 0;
		   board[26][53] <= 0;
		   board[26][54] <= 0;
		   board[26][55] <= 0;
		   board[26][56] <= 0;
		   board[26][57] <= 0;
		   board[26][58] <= 0;
		   board[26][59] <= 0;
		   board[26][60] <= 0;
		   board[26][61] <= 0;
		   board[26][62] <= 0;
		   board[26][63] <= 0;
		   board[27][0] <= 0;
		   board[27][1] <= 0;
		   board[27][2] <= 0;
		   board[27][3] <= 0;
		   board[27][4] <= 0;
		   board[27][5] <= 0;
		   board[27][6] <= 0;
		   board[27][7] <= 0;
		   board[27][8] <= 0;
		   board[27][9] <= 0;
		   board[27][10] <= 0;
		   board[27][11] <= 0;
		   board[27][12] <= 0;
		   board[27][13] <= 0;
		   board[27][14] <= 0;
		   board[27][15] <= 0;
		   board[27][16] <= 0;
		   board[27][17] <= 0;
		   board[27][18] <= 0;
		   board[27][19] <= 0;
		   board[27][20] <= 0;
		   board[27][21] <= 0;
		   board[27][22] <= 0;
		   board[27][23] <= 0;
		   board[27][24] <= 0;
		   board[27][25] <= 0;
		   board[27][26] <= 0;
		   board[27][27] <= 0;
		   board[27][28] <= 0;
		   board[27][29] <= 0;
		   board[27][30] <= 0;
		   board[27][31] <= 0;
		   board[27][32] <= 0;
		   board[27][33] <= 0;
		   board[27][34] <= 0;
		   board[27][35] <= 0;
		   board[27][36] <= 0;
		   board[27][37] <= 0;
		   board[27][38] <= 0;
		   board[27][39] <= 0;
		   board[27][40] <= 0;
		   board[27][41] <= 0;
		   board[27][42] <= 0;
		   board[27][43] <= 0;
		   board[27][44] <= 0;
		   board[27][45] <= 0;
		   board[27][46] <= 0;
		   board[27][47] <= 0;
		   board[27][48] <= 0;
		   board[27][49] <= 0;
		   board[27][50] <= 0;
		   board[27][51] <= 0;
		   board[27][52] <= 0;
		   board[27][53] <= 0;
		   board[27][54] <= 0;
		   board[27][55] <= 0;
		   board[27][56] <= 0;
		   board[27][57] <= 0;
		   board[27][58] <= 0;
		   board[27][59] <= 0;
		   board[27][60] <= 0;
		   board[27][61] <= 0;
		   board[27][62] <= 0;
		   board[27][63] <= 0;
		   board[28][0] <= 0;
		   board[28][1] <= 0;
		   board[28][2] <= 0;
		   board[28][3] <= 0;
		   board[28][4] <= 0;
		   board[28][5] <= 0;
		   board[28][6] <= 0;
		   board[28][7] <= 0;
		   board[28][8] <= 0;
		   board[28][9] <= 0;
		   board[28][10] <= 0;
		   board[28][11] <= 0;
		   board[28][12] <= 0;
		   board[28][13] <= 0;
		   board[28][14] <= 0;
		   board[28][15] <= 0;
		   board[28][16] <= 0;
		   board[28][17] <= 0;
		   board[28][18] <= 0;
		   board[28][19] <= 0;
		   board[28][20] <= 0;
		   board[28][21] <= 0;
		   board[28][22] <= 0;
		   board[28][23] <= 0;
		   board[28][24] <= 0;
		   board[28][25] <= 0;
		   board[28][26] <= 0;
		   board[28][27] <= 0;
		   board[28][28] <= 0;
		   board[28][29] <= 0;
		   board[28][30] <= 0;
		   board[28][31] <= 0;
		   board[28][32] <= 0;
		   board[28][33] <= 0;
		   board[28][34] <= 0;
		   board[28][35] <= 0;
		   board[28][36] <= 0;
		   board[28][37] <= 0;
		   board[28][38] <= 0;
		   board[28][39] <= 0;
		   board[28][40] <= 0;
		   board[28][41] <= 0;
		   board[28][42] <= 0;
		   board[28][43] <= 0;
		   board[28][44] <= 0;
		   board[28][45] <= 0;
		   board[28][46] <= 0;
		   board[28][47] <= 0;
		   board[28][48] <= 0;
		   board[28][49] <= 0;
		   board[28][50] <= 0;
		   board[28][51] <= 0;
		   board[28][52] <= 0;
		   board[28][53] <= 0;
		   board[28][54] <= 0;
		   board[28][55] <= 0;
		   board[28][56] <= 0;
		   board[28][57] <= 0;
		   board[28][58] <= 0;
		   board[28][59] <= 0;
		   board[28][60] <= 0;
		   board[28][61] <= 0;
		   board[28][62] <= 0;
		   board[28][63] <= 0;
		   board[29][0] <= 0;
		   board[29][1] <= 0;
		   board[29][2] <= 0;
		   board[29][3] <= 0;
		   board[29][4] <= 0;
		   board[29][5] <= 0;
		   board[29][6] <= 0;
		   board[29][7] <= 0;
		   board[29][8] <= 0;
		   board[29][9] <= 0;
		   board[29][10] <= 0;
		   board[29][11] <= 0;
		   board[29][12] <= 0;
		   board[29][13] <= 0;
		   board[29][14] <= 0;
		   board[29][15] <= 0;
		   board[29][16] <= 0;
		   board[29][17] <= 0;
		   board[29][18] <= 0;
		   board[29][19] <= 0;
		   board[29][20] <= 0;
		   board[29][21] <= 0;
		   board[29][22] <= 0;
		   board[29][23] <= 0;
		   board[29][24] <= 0;
		   board[29][25] <= 0;
		   board[29][26] <= 0;
		   board[29][27] <= 0;
		   board[29][28] <= 0;
		   board[29][29] <= 0;
		   board[29][30] <= 0;
		   board[29][31] <= 0;
		   board[29][32] <= 0;
		   board[29][33] <= 0;
		   board[29][34] <= 0;
		   board[29][35] <= 0;
		   board[29][36] <= 0;
		   board[29][37] <= 0;
		   board[29][38] <= 0;
		   board[29][39] <= 0;
		   board[29][40] <= 0;
		   board[29][41] <= 0;
		   board[29][42] <= 0;
		   board[29][43] <= 0;
		   board[29][44] <= 0;
		   board[29][45] <= 0;
		   board[29][46] <= 0;
		   board[29][47] <= 0;
		   board[29][48] <= 0;
		   board[29][49] <= 0;
		   board[29][50] <= 0;
		   board[29][51] <= 0;
		   board[29][52] <= 0;
		   board[29][53] <= 0;
		   board[29][54] <= 0;
		   board[29][55] <= 0;
		   board[29][56] <= 0;
		   board[29][57] <= 0;
		   board[29][58] <= 0;
		   board[29][59] <= 0;
		   board[29][60] <= 0;
		   board[29][61] <= 0;
		   board[29][62] <= 0;
		   board[29][63] <= 0;
		   board[30][0] <= 0;
		   board[30][1] <= 0;
		   board[30][2] <= 0;
		   board[30][3] <= 0;
		   board[30][4] <= 0;
		   board[30][5] <= 0;
		   board[30][6] <= 0;
		   board[30][7] <= 0;
		   board[30][8] <= 0;
		   board[30][9] <= 0;
		   board[30][10] <= 0;
		   board[30][11] <= 0;
		   board[30][12] <= 0;
		   board[30][13] <= 0;
		   board[30][14] <= 0;
		   board[30][15] <= 0;
		   board[30][16] <= 0;
		   board[30][17] <= 0;
		   board[30][18] <= 0;
		   board[30][19] <= 0;
		   board[30][20] <= 0;
		   board[30][21] <= 0;
		   board[30][22] <= 0;
		   board[30][23] <= 0;
		   board[30][24] <= 0;
		   board[30][25] <= 0;
		   board[30][26] <= 0;
		   board[30][27] <= 0;
		   board[30][28] <= 0;
		   board[30][29] <= 0;
		   board[30][30] <= 0;
		   board[30][31] <= 0;
		   board[30][32] <= 0;
		   board[30][33] <= 0;
		   board[30][34] <= 0;
		   board[30][35] <= 0;
		   board[30][36] <= 0;
		   board[30][37] <= 0;
		   board[30][38] <= 0;
		   board[30][39] <= 0;
		   board[30][40] <= 0;
		   board[30][41] <= 0;
		   board[30][42] <= 0;
		   board[30][43] <= 0;
		   board[30][44] <= 0;
		   board[30][45] <= 0;
		   board[30][46] <= 0;
		   board[30][47] <= 0;
		   board[30][48] <= 0;
		   board[30][49] <= 0;
		   board[30][50] <= 0;
		   board[30][51] <= 0;
		   board[30][52] <= 0;
		   board[30][53] <= 0;
		   board[30][54] <= 0;
		   board[30][55] <= 0;
		   board[30][56] <= 0;
		   board[30][57] <= 0;
		   board[30][58] <= 0;
		   board[30][59] <= 0;
		   board[30][60] <= 0;
		   board[30][61] <= 0;
		   board[30][62] <= 0;
		   board[30][63] <= 0;
		   board[31][0] <= 0;
		   board[31][1] <= 0;
		   board[31][2] <= 0;
		   board[31][3] <= 0;
		   board[31][4] <= 0;
		   board[31][5] <= 0;
		   board[31][6] <= 0;
		   board[31][7] <= 0;
		   board[31][8] <= 0;
		   board[31][9] <= 0;
		   board[31][10] <= 0;
		   board[31][11] <= 0;
		   board[31][12] <= 0;
		   board[31][13] <= 0;
		   board[31][14] <= 0;
		   board[31][15] <= 0;
		   board[31][16] <= 0;
		   board[31][17] <= 0;
		   board[31][18] <= 0;
		   board[31][19] <= 0;
		   board[31][20] <= 0;
		   board[31][21] <= 0;
		   board[31][22] <= 0;
		   board[31][23] <= 0;
		   board[31][24] <= 0;
		   board[31][25] <= 0;
		   board[31][26] <= 0;
		   board[31][27] <= 0;
		   board[31][28] <= 0;
		   board[31][29] <= 0;
		   board[31][30] <= 0;
		   board[31][31] <= 0;
		   board[31][32] <= 0;
		   board[31][33] <= 0;
		   board[31][34] <= 0;
		   board[31][35] <= 0;
		   board[31][36] <= 0;
		   board[31][37] <= 0;
		   board[31][38] <= 0;
		   board[31][39] <= 0;
		   board[31][40] <= 0;
		   board[31][41] <= 0;
		   board[31][42] <= 0;
		   board[31][43] <= 0;
		   board[31][44] <= 0;
		   board[31][45] <= 0;
		   board[31][46] <= 0;
		   board[31][47] <= 0;
		   board[31][48] <= 0;
		   board[31][49] <= 0;
		   board[31][50] <= 0;
		   board[31][51] <= 0;
		   board[31][52] <= 0;
		   board[31][53] <= 0;
		   board[31][54] <= 0;
		   board[31][55] <= 0;
		   board[31][56] <= 0;
		   board[31][57] <= 0;
		   board[31][58] <= 0;
		   board[31][59] <= 0;
		   board[31][60] <= 0;
		   board[31][61] <= 0;
		   board[31][62] <= 0;
		   board[31][63] <= 0;
		   board[32][0] <= 0;
		   board[32][1] <= 0;
		   board[32][2] <= 0;
		   board[32][3] <= 0;
		   board[32][4] <= 0;
		   board[32][5] <= 0;
		   board[32][6] <= 0;
		   board[32][7] <= 0;
		   board[32][8] <= 0;
		   board[32][9] <= 0;
		   board[32][10] <= 0;
		   board[32][11] <= 0;
		   board[32][12] <= 0;
		   board[32][13] <= 0;
		   board[32][14] <= 0;
		   board[32][15] <= 0;
		   board[32][16] <= 0;
		   board[32][17] <= 0;
		   board[32][18] <= 0;
		   board[32][19] <= 0;
		   board[32][20] <= 0;
		   board[32][21] <= 0;
		   board[32][22] <= 0;
		   board[32][23] <= 0;
		   board[32][24] <= 0;
		   board[32][25] <= 0;
		   board[32][26] <= 0;
		   board[32][27] <= 0;
		   board[32][28] <= 0;
		   board[32][29] <= 0;
		   board[32][30] <= 0;
		   board[32][31] <= 0;
		   board[32][32] <= 0;
		   board[32][33] <= 0;
		   board[32][34] <= 0;
		   board[32][35] <= 0;
		   board[32][36] <= 0;
		   board[32][37] <= 0;
		   board[32][38] <= 0;
		   board[32][39] <= 0;
		   board[32][40] <= 0;
		   board[32][41] <= 0;
		   board[32][42] <= 0;
		   board[32][43] <= 0;
		   board[32][44] <= 0;
		   board[32][45] <= 0;
		   board[32][46] <= 0;
		   board[32][47] <= 0;
		   board[32][48] <= 0;
		   board[32][49] <= 0;
		   board[32][50] <= 0;
		   board[32][51] <= 0;
		   board[32][52] <= 0;
		   board[32][53] <= 0;
		   board[32][54] <= 0;
		   board[32][55] <= 0;
		   board[32][56] <= 0;
		   board[32][57] <= 0;
		   board[32][58] <= 0;
		   board[32][59] <= 0;
		   board[32][60] <= 0;
		   board[32][61] <= 0;
		   board[32][62] <= 0;
		   board[32][63] <= 0;
		   board[33][0] <= 0;
		   board[33][1] <= 0;
		   board[33][2] <= 0;
		   board[33][3] <= 0;
		   board[33][4] <= 0;
		   board[33][5] <= 0;
		   board[33][6] <= 0;
		   board[33][7] <= 0;
		   board[33][8] <= 0;
		   board[33][9] <= 0;
		   board[33][10] <= 0;
		   board[33][11] <= 0;
		   board[33][12] <= 0;
		   board[33][13] <= 0;
		   board[33][14] <= 0;
		   board[33][15] <= 0;
		   board[33][16] <= 0;
		   board[33][17] <= 0;
		   board[33][18] <= 0;
		   board[33][19] <= 0;
		   board[33][20] <= 0;
		   board[33][21] <= 0;
		   board[33][22] <= 0;
		   board[33][23] <= 0;
		   board[33][24] <= 0;
		   board[33][25] <= 0;
		   board[33][26] <= 0;
		   board[33][27] <= 0;
		   board[33][28] <= 0;
		   board[33][29] <= 0;
		   board[33][30] <= 0;
		   board[33][31] <= 0;
		   board[33][32] <= 0;
		   board[33][33] <= 0;
		   board[33][34] <= 0;
		   board[33][35] <= 0;
		   board[33][36] <= 0;
		   board[33][37] <= 0;
		   board[33][38] <= 0;
		   board[33][39] <= 0;
		   board[33][40] <= 0;
		   board[33][41] <= 0;
		   board[33][42] <= 0;
		   board[33][43] <= 0;
		   board[33][44] <= 0;
		   board[33][45] <= 0;
		   board[33][46] <= 0;
		   board[33][47] <= 0;
		   board[33][48] <= 0;
		   board[33][49] <= 0;
		   board[33][50] <= 0;
		   board[33][51] <= 0;
		   board[33][52] <= 0;
		   board[33][53] <= 0;
		   board[33][54] <= 0;
		   board[33][55] <= 0;
		   board[33][56] <= 0;
		   board[33][57] <= 0;
		   board[33][58] <= 0;
		   board[33][59] <= 0;
		   board[33][60] <= 0;
		   board[33][61] <= 0;
		   board[33][62] <= 0;
		   board[33][63] <= 0;
		   board[34][0] <= 0;
		   board[34][1] <= 0;
		   board[34][2] <= 0;
		   board[34][3] <= 0;
		   board[34][4] <= 0;
		   board[34][5] <= 0;
		   board[34][6] <= 0;
		   board[34][7] <= 0;
		   board[34][8] <= 0;
		   board[34][9] <= 0;
		   board[34][10] <= 0;
		   board[34][11] <= 0;
		   board[34][12] <= 0;
		   board[34][13] <= 0;
		   board[34][14] <= 0;
		   board[34][15] <= 0;
		   board[34][16] <= 0;
		   board[34][17] <= 0;
		   board[34][18] <= 0;
		   board[34][19] <= 0;
		   board[34][20] <= 0;
		   board[34][21] <= 0;
		   board[34][22] <= 0;
		   board[34][23] <= 0;
		   board[34][24] <= 0;
		   board[34][25] <= 0;
		   board[34][26] <= 0;
		   board[34][27] <= 0;
		   board[34][28] <= 0;
		   board[34][29] <= 0;
		   board[34][30] <= 0;
		   board[34][31] <= 0;
		   board[34][32] <= 0;
		   board[34][33] <= 0;
		   board[34][34] <= 0;
		   board[34][35] <= 0;
		   board[34][36] <= 0;
		   board[34][37] <= 0;
		   board[34][38] <= 0;
		   board[34][39] <= 0;
		   board[34][40] <= 0;
		   board[34][41] <= 0;
		   board[34][42] <= 0;
		   board[34][43] <= 0;
		   board[34][44] <= 0;
		   board[34][45] <= 0;
		   board[34][46] <= 0;
		   board[34][47] <= 0;
		   board[34][48] <= 0;
		   board[34][49] <= 0;
		   board[34][50] <= 0;
		   board[34][51] <= 0;
		   board[34][52] <= 0;
		   board[34][53] <= 0;
		   board[34][54] <= 0;
		   board[34][55] <= 0;
		   board[34][56] <= 0;
		   board[34][57] <= 0;
		   board[34][58] <= 0;
		   board[34][59] <= 0;
		   board[34][60] <= 0;
		   board[34][61] <= 0;
		   board[34][62] <= 0;
		   board[34][63] <= 0;
		   board[35][0] <= 0;
		   board[35][1] <= 0;
		   board[35][2] <= 0;
		   board[35][3] <= 0;
		   board[35][4] <= 0;
		   board[35][5] <= 0;
		   board[35][6] <= 0;
		   board[35][7] <= 0;
		   board[35][8] <= 0;
		   board[35][9] <= 0;
		   board[35][10] <= 0;
		   board[35][11] <= 0;
		   board[35][12] <= 0;
		   board[35][13] <= 0;
		   board[35][14] <= 0;
		   board[35][15] <= 0;
		   board[35][16] <= 0;
		   board[35][17] <= 0;
		   board[35][18] <= 0;
		   board[35][19] <= 0;
		   board[35][20] <= 0;
		   board[35][21] <= 0;
		   board[35][22] <= 0;
		   board[35][23] <= 0;
		   board[35][24] <= 0;
		   board[35][25] <= 0;
		   board[35][26] <= 0;
		   board[35][27] <= 0;
		   board[35][28] <= 0;
		   board[35][29] <= 0;
		   board[35][30] <= 0;
		   board[35][31] <= 0;
		   board[35][32] <= 0;
		   board[35][33] <= 0;
		   board[35][34] <= 0;
		   board[35][35] <= 0;
		   board[35][36] <= 0;
		   board[35][37] <= 0;
		   board[35][38] <= 0;
		   board[35][39] <= 0;
		   board[35][40] <= 0;
		   board[35][41] <= 0;
		   board[35][42] <= 0;
		   board[35][43] <= 0;
		   board[35][44] <= 0;
		   board[35][45] <= 0;
		   board[35][46] <= 0;
		   board[35][47] <= 0;
		   board[35][48] <= 0;
		   board[35][49] <= 0;
		   board[35][50] <= 0;
		   board[35][51] <= 0;
		   board[35][52] <= 0;
		   board[35][53] <= 0;
		   board[35][54] <= 0;
		   board[35][55] <= 0;
		   board[35][56] <= 0;
		   board[35][57] <= 0;
		   board[35][58] <= 0;
		   board[35][59] <= 0;
		   board[35][60] <= 0;
		   board[35][61] <= 0;
		   board[35][62] <= 0;
		   board[35][63] <= 0;
		   board[36][0] <= 0;
		   board[36][1] <= 0;
		   board[36][2] <= 0;
		   board[36][3] <= 0;
		   board[36][4] <= 0;
		   board[36][5] <= 0;
		   board[36][6] <= 0;
		   board[36][7] <= 0;
		   board[36][8] <= 0;
		   board[36][9] <= 0;
		   board[36][10] <= 0;
		   board[36][11] <= 0;
		   board[36][12] <= 0;
		   board[36][13] <= 0;
		   board[36][14] <= 0;
		   board[36][15] <= 0;
		   board[36][16] <= 0;
		   board[36][17] <= 0;
		   board[36][18] <= 0;
		   board[36][19] <= 0;
		   board[36][20] <= 0;
		   board[36][21] <= 0;
		   board[36][22] <= 0;
		   board[36][23] <= 0;
		   board[36][24] <= 0;
		   board[36][25] <= 0;
		   board[36][26] <= 0;
		   board[36][27] <= 0;
		   board[36][28] <= 0;
		   board[36][29] <= 0;
		   board[36][30] <= 0;
		   board[36][31] <= 0;
		   board[36][32] <= 0;
		   board[36][33] <= 0;
		   board[36][34] <= 0;
		   board[36][35] <= 0;
		   board[36][36] <= 0;
		   board[36][37] <= 0;
		   board[36][38] <= 0;
		   board[36][39] <= 0;
		   board[36][40] <= 0;
		   board[36][41] <= 0;
		   board[36][42] <= 0;
		   board[36][43] <= 0;
		   board[36][44] <= 0;
		   board[36][45] <= 0;
		   board[36][46] <= 0;
		   board[36][47] <= 0;
		   board[36][48] <= 0;
		   board[36][49] <= 0;
		   board[36][50] <= 0;
		   board[36][51] <= 0;
		   board[36][52] <= 0;
		   board[36][53] <= 0;
		   board[36][54] <= 0;
		   board[36][55] <= 0;
		   board[36][56] <= 0;
		   board[36][57] <= 0;
		   board[36][58] <= 0;
		   board[36][59] <= 0;
		   board[36][60] <= 0;
		   board[36][61] <= 0;
		   board[36][62] <= 0;
		   board[36][63] <= 0;
		   board[37][0] <= 0;
		   board[37][1] <= 0;
		   board[37][2] <= 0;
		   board[37][3] <= 0;
		   board[37][4] <= 0;
		   board[37][5] <= 0;
		   board[37][6] <= 0;
		   board[37][7] <= 0;
		   board[37][8] <= 0;
		   board[37][9] <= 0;
		   board[37][10] <= 0;
		   board[37][11] <= 0;
		   board[37][12] <= 0;
		   board[37][13] <= 0;
		   board[37][14] <= 0;
		   board[37][15] <= 0;
		   board[37][16] <= 0;
		   board[37][17] <= 0;
		   board[37][18] <= 0;
		   board[37][19] <= 0;
		   board[37][20] <= 0;
		   board[37][21] <= 0;
		   board[37][22] <= 0;
		   board[37][23] <= 0;
		   board[37][24] <= 0;
		   board[37][25] <= 0;
		   board[37][26] <= 0;
		   board[37][27] <= 0;
		   board[37][28] <= 0;
		   board[37][29] <= 0;
		   board[37][30] <= 0;
		   board[37][31] <= 0;
		   board[37][32] <= 0;
		   board[37][33] <= 0;
		   board[37][34] <= 0;
		   board[37][35] <= 0;
		   board[37][36] <= 0;
		   board[37][37] <= 0;
		   board[37][38] <= 0;
		   board[37][39] <= 0;
		   board[37][40] <= 0;
		   board[37][41] <= 0;
		   board[37][42] <= 0;
		   board[37][43] <= 0;
		   board[37][44] <= 0;
		   board[37][45] <= 0;
		   board[37][46] <= 0;
		   board[37][47] <= 0;
		   board[37][48] <= 0;
		   board[37][49] <= 0;
		   board[37][50] <= 0;
		   board[37][51] <= 0;
		   board[37][52] <= 0;
		   board[37][53] <= 0;
		   board[37][54] <= 0;
		   board[37][55] <= 0;
		   board[37][56] <= 0;
		   board[37][57] <= 0;
		   board[37][58] <= 0;
		   board[37][59] <= 0;
		   board[37][60] <= 0;
		   board[37][61] <= 0;
		   board[37][62] <= 0;
		   board[37][63] <= 0;
		   board[38][0] <= 0;
		   board[38][1] <= 0;
		   board[38][2] <= 0;
		   board[38][3] <= 0;
		   board[38][4] <= 0;
		   board[38][5] <= 0;
		   board[38][6] <= 0;
		   board[38][7] <= 0;
		   board[38][8] <= 0;
		   board[38][9] <= 0;
		   board[38][10] <= 0;
		   board[38][11] <= 0;
		   board[38][12] <= 0;
		   board[38][13] <= 0;
		   board[38][14] <= 0;
		   board[38][15] <= 0;
		   board[38][16] <= 0;
		   board[38][17] <= 0;
		   board[38][18] <= 0;
		   board[38][19] <= 0;
		   board[38][20] <= 0;
		   board[38][21] <= 0;
		   board[38][22] <= 0;
		   board[38][23] <= 0;
		   board[38][24] <= 0;
		   board[38][25] <= 0;
		   board[38][26] <= 0;
		   board[38][27] <= 0;
		   board[38][28] <= 0;
		   board[38][29] <= 0;
		   board[38][30] <= 0;
		   board[38][31] <= 0;
		   board[38][32] <= 0;
		   board[38][33] <= 0;
		   board[38][34] <= 0;
		   board[38][35] <= 0;
		   board[38][36] <= 0;
		   board[38][37] <= 0;
		   board[38][38] <= 0;
		   board[38][39] <= 0;
		   board[38][40] <= 0;
		   board[38][41] <= 0;
		   board[38][42] <= 0;
		   board[38][43] <= 0;
		   board[38][44] <= 0;
		   board[38][45] <= 0;
		   board[38][46] <= 0;
		   board[38][47] <= 0;
		   board[38][48] <= 0;
		   board[38][49] <= 0;
		   board[38][50] <= 0;
		   board[38][51] <= 0;
		   board[38][52] <= 0;
		   board[38][53] <= 0;
		   board[38][54] <= 0;
		   board[38][55] <= 0;
		   board[38][56] <= 0;
		   board[38][57] <= 0;
		   board[38][58] <= 0;
		   board[38][59] <= 0;
		   board[38][60] <= 0;
		   board[38][61] <= 0;
		   board[38][62] <= 0;
		   board[38][63] <= 0;
		   board[39][0] <= 0;
		   board[39][1] <= 0;
		   board[39][2] <= 0;
		   board[39][3] <= 0;
		   board[39][4] <= 0;
		   board[39][5] <= 0;
		   board[39][6] <= 0;
		   board[39][7] <= 0;
		   board[39][8] <= 0;
		   board[39][9] <= 0;
		   board[39][10] <= 0;
		   board[39][11] <= 0;
		   board[39][12] <= 0;
		   board[39][13] <= 0;
		   board[39][14] <= 0;
		   board[39][15] <= 0;
		   board[39][16] <= 0;
		   board[39][17] <= 0;
		   board[39][18] <= 0;
		   board[39][19] <= 0;
		   board[39][20] <= 0;
		   board[39][21] <= 0;
		   board[39][22] <= 0;
		   board[39][23] <= 0;
		   board[39][24] <= 0;
		   board[39][25] <= 0;
		   board[39][26] <= 0;
		   board[39][27] <= 0;
		   board[39][28] <= 0;
		   board[39][29] <= 0;
		   board[39][30] <= 0;
		   board[39][31] <= 0;
		   board[39][32] <= 0;
		   board[39][33] <= 0;
		   board[39][34] <= 0;
		   board[39][35] <= 0;
		   board[39][36] <= 0;
		   board[39][37] <= 0;
		   board[39][38] <= 0;
		   board[39][39] <= 0;
		   board[39][40] <= 0;
		   board[39][41] <= 0;
		   board[39][42] <= 0;
		   board[39][43] <= 0;
		   board[39][44] <= 0;
		   board[39][45] <= 0;
		   board[39][46] <= 0;
		   board[39][47] <= 0;
		   board[39][48] <= 0;
		   board[39][49] <= 0;
		   board[39][50] <= 0;
		   board[39][51] <= 0;
		   board[39][52] <= 0;
		   board[39][53] <= 0;
		   board[39][54] <= 0;
		   board[39][55] <= 0;
		   board[39][56] <= 0;
		   board[39][57] <= 0;
		   board[39][58] <= 0;
		   board[39][59] <= 0;
		   board[39][60] <= 0;
		   board[39][61] <= 0;
		   board[39][62] <= 0;
		   board[39][63] <= 0;
		   board[40][0] <= 0;
		   board[40][1] <= 0;
		   board[40][2] <= 0;
		   board[40][3] <= 0;
		   board[40][4] <= 0;
		   board[40][5] <= 0;
		   board[40][6] <= 0;
		   board[40][7] <= 0;
		   board[40][8] <= 0;
		   board[40][9] <= 0;
		   board[40][10] <= 0;
		   board[40][11] <= 0;
		   board[40][12] <= 0;
		   board[40][13] <= 0;
		   board[40][14] <= 0;
		   board[40][15] <= 0;
		   board[40][16] <= 0;
		   board[40][17] <= 0;
		   board[40][18] <= 0;
		   board[40][19] <= 0;
		   board[40][20] <= 0;
		   board[40][21] <= 0;
		   board[40][22] <= 0;
		   board[40][23] <= 0;
		   board[40][24] <= 0;
		   board[40][25] <= 0;
		   board[40][26] <= 0;
		   board[40][27] <= 0;
		   board[40][28] <= 0;
		   board[40][29] <= 0;
		   board[40][30] <= 0;
		   board[40][31] <= 0;
		   board[40][32] <= 0;
		   board[40][33] <= 0;
		   board[40][34] <= 0;
		   board[40][35] <= 0;
		   board[40][36] <= 0;
		   board[40][37] <= 0;
		   board[40][38] <= 0;
		   board[40][39] <= 0;
		   board[40][40] <= 0;
		   board[40][41] <= 0;
		   board[40][42] <= 0;
		   board[40][43] <= 0;
		   board[40][44] <= 0;
		   board[40][45] <= 0;
		   board[40][46] <= 0;
		   board[40][47] <= 0;
		   board[40][48] <= 0;
		   board[40][49] <= 0;
		   board[40][50] <= 0;
		   board[40][51] <= 0;
		   board[40][52] <= 0;
		   board[40][53] <= 0;
		   board[40][54] <= 0;
		   board[40][55] <= 0;
		   board[40][56] <= 0;
		   board[40][57] <= 0;
		   board[40][58] <= 0;
		   board[40][59] <= 0;
		   board[40][60] <= 0;
		   board[40][61] <= 0;
		   board[40][62] <= 0;
		   board[40][63] <= 0;
		   board[41][0] <= 0;
		   board[41][1] <= 0;
		   board[41][2] <= 0;
		   board[41][3] <= 0;
		   board[41][4] <= 0;
		   board[41][5] <= 0;
		   board[41][6] <= 0;
		   board[41][7] <= 0;
		   board[41][8] <= 0;
		   board[41][9] <= 0;
		   board[41][10] <= 0;
		   board[41][11] <= 0;
		   board[41][12] <= 0;
		   board[41][13] <= 0;
		   board[41][14] <= 0;
		   board[41][15] <= 0;
		   board[41][16] <= 0;
		   board[41][17] <= 0;
		   board[41][18] <= 0;
		   board[41][19] <= 0;
		   board[41][20] <= 0;
		   board[41][21] <= 0;
		   board[41][22] <= 0;
		   board[41][23] <= 0;
		   board[41][24] <= 0;
		   board[41][25] <= 0;
		   board[41][26] <= 0;
		   board[41][27] <= 0;
		   board[41][28] <= 0;
		   board[41][29] <= 0;
		   board[41][30] <= 0;
		   board[41][31] <= 0;
		   board[41][32] <= 0;
		   board[41][33] <= 0;
		   board[41][34] <= 0;
		   board[41][35] <= 0;
		   board[41][36] <= 0;
		   board[41][37] <= 0;
		   board[41][38] <= 0;
		   board[41][39] <= 0;
		   board[41][40] <= 0;
		   board[41][41] <= 0;
		   board[41][42] <= 0;
		   board[41][43] <= 0;
		   board[41][44] <= 0;
		   board[41][45] <= 0;
		   board[41][46] <= 0;
		   board[41][47] <= 0;
		   board[41][48] <= 0;
		   board[41][49] <= 0;
		   board[41][50] <= 0;
		   board[41][51] <= 0;
		   board[41][52] <= 0;
		   board[41][53] <= 0;
		   board[41][54] <= 0;
		   board[41][55] <= 0;
		   board[41][56] <= 0;
		   board[41][57] <= 0;
		   board[41][58] <= 0;
		   board[41][59] <= 0;
		   board[41][60] <= 0;
		   board[41][61] <= 0;
		   board[41][62] <= 0;
		   board[41][63] <= 0;
		   board[42][0] <= 0;
		   board[42][1] <= 0;
		   board[42][2] <= 0;
		   board[42][3] <= 0;
		   board[42][4] <= 0;
		   board[42][5] <= 0;
		   board[42][6] <= 0;
		   board[42][7] <= 0;
		   board[42][8] <= 0;
		   board[42][9] <= 0;
		   board[42][10] <= 0;
		   board[42][11] <= 0;
		   board[42][12] <= 0;
		   board[42][13] <= 0;
		   board[42][14] <= 0;
		   board[42][15] <= 0;
		   board[42][16] <= 0;
		   board[42][17] <= 0;
		   board[42][18] <= 0;
		   board[42][19] <= 0;
		   board[42][20] <= 0;
		   board[42][21] <= 0;
		   board[42][22] <= 0;
		   board[42][23] <= 0;
		   board[42][24] <= 0;
		   board[42][25] <= 0;
		   board[42][26] <= 0;
		   board[42][27] <= 0;
		   board[42][28] <= 0;
		   board[42][29] <= 0;
		   board[42][30] <= 0;
		   board[42][31] <= 0;
		   board[42][32] <= 0;
		   board[42][33] <= 0;
		   board[42][34] <= 0;
		   board[42][35] <= 0;
		   board[42][36] <= 0;
		   board[42][37] <= 0;
		   board[42][38] <= 0;
		   board[42][39] <= 0;
		   board[42][40] <= 0;
		   board[42][41] <= 0;
		   board[42][42] <= 0;
		   board[42][43] <= 0;
		   board[42][44] <= 0;
		   board[42][45] <= 0;
		   board[42][46] <= 0;
		   board[42][47] <= 0;
		   board[42][48] <= 0;
		   board[42][49] <= 0;
		   board[42][50] <= 0;
		   board[42][51] <= 0;
		   board[42][52] <= 0;
		   board[42][53] <= 0;
		   board[42][54] <= 0;
		   board[42][55] <= 0;
		   board[42][56] <= 0;
		   board[42][57] <= 0;
		   board[42][58] <= 0;
		   board[42][59] <= 0;
		   board[42][60] <= 0;
		   board[42][61] <= 0;
		   board[42][62] <= 0;
		   board[42][63] <= 0;
		   board[43][0] <= 0;
		   board[43][1] <= 0;
		   board[43][2] <= 0;
		   board[43][3] <= 0;
		   board[43][4] <= 0;
		   board[43][5] <= 0;
		   board[43][6] <= 0;
		   board[43][7] <= 0;
		   board[43][8] <= 0;
		   board[43][9] <= 0;
		   board[43][10] <= 0;
		   board[43][11] <= 0;
		   board[43][12] <= 0;
		   board[43][13] <= 0;
		   board[43][14] <= 0;
		   board[43][15] <= 0;
		   board[43][16] <= 0;
		   board[43][17] <= 0;
		   board[43][18] <= 0;
		   board[43][19] <= 0;
		   board[43][20] <= 0;
		   board[43][21] <= 0;
		   board[43][22] <= 0;
		   board[43][23] <= 0;
		   board[43][24] <= 0;
		   board[43][25] <= 0;
		   board[43][26] <= 0;
		   board[43][27] <= 0;
		   board[43][28] <= 0;
		   board[43][29] <= 0;
		   board[43][30] <= 0;
		   board[43][31] <= 0;
		   board[43][32] <= 0;
		   board[43][33] <= 0;
		   board[43][34] <= 0;
		   board[43][35] <= 0;
		   board[43][36] <= 0;
		   board[43][37] <= 0;
		   board[43][38] <= 0;
		   board[43][39] <= 0;
		   board[43][40] <= 0;
		   board[43][41] <= 0;
		   board[43][42] <= 0;
		   board[43][43] <= 0;
		   board[43][44] <= 0;
		   board[43][45] <= 0;
		   board[43][46] <= 0;
		   board[43][47] <= 0;
		   board[43][48] <= 0;
		   board[43][49] <= 0;
		   board[43][50] <= 0;
		   board[43][51] <= 0;
		   board[43][52] <= 0;
		   board[43][53] <= 0;
		   board[43][54] <= 0;
		   board[43][55] <= 0;
		   board[43][56] <= 0;
		   board[43][57] <= 0;
		   board[43][58] <= 0;
		   board[43][59] <= 0;
		   board[43][60] <= 0;
		   board[43][61] <= 0;
		   board[43][62] <= 0;
		   board[43][63] <= 0;
		   board[44][0] <= 0;
		   board[44][1] <= 0;
		   board[44][2] <= 0;
		   board[44][3] <= 0;
		   board[44][4] <= 0;
		   board[44][5] <= 0;
		   board[44][6] <= 0;
		   board[44][7] <= 0;
		   board[44][8] <= 0;
		   board[44][9] <= 0;
		   board[44][10] <= 0;
		   board[44][11] <= 0;
		   board[44][12] <= 0;
		   board[44][13] <= 0;
		   board[44][14] <= 0;
		   board[44][15] <= 0;
		   board[44][16] <= 0;
		   board[44][17] <= 0;
		   board[44][18] <= 0;
		   board[44][19] <= 0;
		   board[44][20] <= 0;
		   board[44][21] <= 0;
		   board[44][22] <= 0;
		   board[44][23] <= 0;
		   board[44][24] <= 0;
		   board[44][25] <= 0;
		   board[44][26] <= 0;
		   board[44][27] <= 0;
		   board[44][28] <= 0;
		   board[44][29] <= 0;
		   board[44][30] <= 0;
		   board[44][31] <= 0;
		   board[44][32] <= 0;
		   board[44][33] <= 0;
		   board[44][34] <= 0;
		   board[44][35] <= 0;
		   board[44][36] <= 0;
		   board[44][37] <= 0;
		   board[44][38] <= 0;
		   board[44][39] <= 0;
		   board[44][40] <= 0;
		   board[44][41] <= 0;
		   board[44][42] <= 0;
		   board[44][43] <= 0;
		   board[44][44] <= 0;
		   board[44][45] <= 0;
		   board[44][46] <= 0;
		   board[44][47] <= 0;
		   board[44][48] <= 0;
		   board[44][49] <= 0;
		   board[44][50] <= 0;
		   board[44][51] <= 0;
		   board[44][52] <= 0;
		   board[44][53] <= 0;
		   board[44][54] <= 0;
		   board[44][55] <= 0;
		   board[44][56] <= 0;
		   board[44][57] <= 0;
		   board[44][58] <= 0;
		   board[44][59] <= 0;
		   board[44][60] <= 0;
		   board[44][61] <= 0;
		   board[44][62] <= 0;
		   board[44][63] <= 0;
		   board[45][0] <= 0;
		   board[45][1] <= 0;
		   board[45][2] <= 0;
		   board[45][3] <= 0;
		   board[45][4] <= 0;
		   board[45][5] <= 0;
		   board[45][6] <= 0;
		   board[45][7] <= 0;
		   board[45][8] <= 0;
		   board[45][9] <= 0;
		   board[45][10] <= 0;
		   board[45][11] <= 0;
		   board[45][12] <= 0;
		   board[45][13] <= 0;
		   board[45][14] <= 0;
		   board[45][15] <= 0;
		   board[45][16] <= 0;
		   board[45][17] <= 0;
		   board[45][18] <= 0;
		   board[45][19] <= 0;
		   board[45][20] <= 0;
		   board[45][21] <= 0;
		   board[45][22] <= 0;
		   board[45][23] <= 0;
		   board[45][24] <= 0;
		   board[45][25] <= 0;
		   board[45][26] <= 0;
		   board[45][27] <= 0;
		   board[45][28] <= 0;
		   board[45][29] <= 0;
		   board[45][30] <= 0;
		   board[45][31] <= 0;
		   board[45][32] <= 0;
		   board[45][33] <= 0;
		   board[45][34] <= 0;
		   board[45][35] <= 0;
		   board[45][36] <= 0;
		   board[45][37] <= 0;
		   board[45][38] <= 0;
		   board[45][39] <= 0;
		   board[45][40] <= 0;
		   board[45][41] <= 0;
		   board[45][42] <= 0;
		   board[45][43] <= 0;
		   board[45][44] <= 0;
		   board[45][45] <= 0;
		   board[45][46] <= 0;
		   board[45][47] <= 0;
		   board[45][48] <= 0;
		   board[45][49] <= 0;
		   board[45][50] <= 0;
		   board[45][51] <= 0;
		   board[45][52] <= 0;
		   board[45][53] <= 0;
		   board[45][54] <= 0;
		   board[45][55] <= 0;
		   board[45][56] <= 0;
		   board[45][57] <= 0;
		   board[45][58] <= 0;
		   board[45][59] <= 0;
		   board[45][60] <= 0;
		   board[45][61] <= 0;
		   board[45][62] <= 0;
		   board[45][63] <= 0;
		   board[46][0] <= 0;
		   board[46][1] <= 0;
		   board[46][2] <= 0;
		   board[46][3] <= 0;
		   board[46][4] <= 0;
		   board[46][5] <= 0;
		   board[46][6] <= 0;
		   board[46][7] <= 0;
		   board[46][8] <= 0;
		   board[46][9] <= 0;
		   board[46][10] <= 0;
		   board[46][11] <= 0;
		   board[46][12] <= 0;
		   board[46][13] <= 0;
		   board[46][14] <= 0;
		   board[46][15] <= 0;
		   board[46][16] <= 0;
		   board[46][17] <= 0;
		   board[46][18] <= 0;
		   board[46][19] <= 0;
		   board[46][20] <= 0;
		   board[46][21] <= 0;
		   board[46][22] <= 0;
		   board[46][23] <= 0;
		   board[46][24] <= 0;
		   board[46][25] <= 0;
		   board[46][26] <= 0;
		   board[46][27] <= 0;
		   board[46][28] <= 0;
		   board[46][29] <= 0;
		   board[46][30] <= 0;
		   board[46][31] <= 0;
		   board[46][32] <= 0;
		   board[46][33] <= 0;
		   board[46][34] <= 0;
		   board[46][35] <= 0;
		   board[46][36] <= 0;
		   board[46][37] <= 0;
		   board[46][38] <= 0;
		   board[46][39] <= 0;
		   board[46][40] <= 0;
		   board[46][41] <= 0;
		   board[46][42] <= 0;
		   board[46][43] <= 0;
		   board[46][44] <= 0;
		   board[46][45] <= 0;
		   board[46][46] <= 0;
		   board[46][47] <= 0;
		   board[46][48] <= 0;
		   board[46][49] <= 0;
		   board[46][50] <= 0;
		   board[46][51] <= 0;
		   board[46][52] <= 0;
		   board[46][53] <= 0;
		   board[46][54] <= 0;
		   board[46][55] <= 0;
		   board[46][56] <= 0;
		   board[46][57] <= 0;
		   board[46][58] <= 0;
		   board[46][59] <= 0;
		   board[46][60] <= 0;
		   board[46][61] <= 0;
		   board[46][62] <= 0;
		   board[46][63] <= 0;
		   board[47][0] <= 0;
		   board[47][1] <= 0;
		   board[47][2] <= 0;
		   board[47][3] <= 0;
		   board[47][4] <= 0;
		   board[47][5] <= 0;
		   board[47][6] <= 0;
		   board[47][7] <= 0;
		   board[47][8] <= 0;
		   board[47][9] <= 0;
		   board[47][10] <= 0;
		   board[47][11] <= 0;
		   board[47][12] <= 0;
		   board[47][13] <= 0;
		   board[47][14] <= 0;
		   board[47][15] <= 0;
		   board[47][16] <= 0;
		   board[47][17] <= 0;
		   board[47][18] <= 0;
		   board[47][19] <= 0;
		   board[47][20] <= 0;
		   board[47][21] <= 0;
		   board[47][22] <= 0;
		   board[47][23] <= 0;
		   board[47][24] <= 0;
		   board[47][25] <= 0;
		   board[47][26] <= 0;
		   board[47][27] <= 0;
		   board[47][28] <= 0;
		   board[47][29] <= 0;
		   board[47][30] <= 0;
		   board[47][31] <= 0;
		   board[47][32] <= 0;
		   board[47][33] <= 0;
		   board[47][34] <= 0;
		   board[47][35] <= 0;
		   board[47][36] <= 0;
		   board[47][37] <= 0;
		   board[47][38] <= 0;
		   board[47][39] <= 0;
		   board[47][40] <= 0;
		   board[47][41] <= 0;
		   board[47][42] <= 0;
		   board[47][43] <= 0;
		   board[47][44] <= 0;
		   board[47][45] <= 0;
		   board[47][46] <= 0;
		   board[47][47] <= 0;
		   board[47][48] <= 0;
		   board[47][49] <= 0;
		   board[47][50] <= 0;
		   board[47][51] <= 0;
		   board[47][52] <= 0;
		   board[47][53] <= 0;
		   board[47][54] <= 0;
		   board[47][55] <= 0;
		   board[47][56] <= 0;
		   board[47][57] <= 0;
		   board[47][58] <= 0;
		   board[47][59] <= 0;
		   board[47][60] <= 0;
		   board[47][61] <= 0;
		   board[47][62] <= 0;
		   board[47][63] <= 0;
		end else begin
			for (i = 0; i < ROWS; i = i + 1) begin
				for (j = 0; j < COLUMNS; j = j + 1) begin
					board[i][j] <= next_board[i][j];
				end
			end
		end
	end
	
	always @(*) begin
		integer i, j, neighbors;
		
		for (i = 1; i < ROWS - 1; i = i + 1) begin
			for (j = 1; j < COLUMNS - 1; j = j + 1) begin
				neighbors = board[i-1][j-1] + board[i][j-1] + board[i+1][j-1] +
								board[i-1][j]   +                 board[i+1][j]   +
								board[i-1][j+1] + board[i][j+1] + board[i+1][j+1];
								
				if (board[i][j]) begin
					next_board[i][j] = neighbors == 2 || neighbors == 3;
				end else begin
					next_board[i][j] = neighbors == 3;
				end
			end
		end
	end
	
	assign pixel = board[row][column];
endmodule